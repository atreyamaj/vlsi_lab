magic
tech scmos
timestamp 1199203464
<< ab >>
rect 0 0 64 72
<< nwell >>
rect -5 32 69 77
<< pwell >>
rect -5 -5 69 32
<< poly >>
rect 11 67 34 69
rect 11 61 13 67
rect 9 58 13 61
rect 22 59 24 63
rect 32 59 34 67
rect 42 65 44 70
rect 49 65 51 70
rect 9 55 11 58
rect 22 44 24 47
rect 9 40 11 43
rect 22 42 27 44
rect 32 42 34 47
rect 42 42 44 47
rect 49 44 51 47
rect 9 38 15 40
rect 9 36 11 38
rect 13 36 15 38
rect 9 34 15 36
rect 13 31 15 34
rect 25 35 27 42
rect 39 40 44 42
rect 48 42 54 44
rect 48 40 50 42
rect 52 40 54 42
rect 25 33 31 35
rect 25 31 27 33
rect 29 31 31 33
rect 13 29 19 31
rect 25 29 31 31
rect 17 26 19 29
rect 29 26 31 29
rect 39 26 41 40
rect 48 38 54 40
rect 49 26 51 38
rect 7 16 13 18
rect 7 14 9 16
rect 11 14 13 16
rect 17 15 19 20
rect 7 12 13 14
rect 29 15 31 20
rect 11 10 13 12
rect 39 10 41 20
rect 49 15 51 20
rect 55 16 61 18
rect 55 14 57 16
rect 59 14 61 16
rect 55 12 61 14
rect 55 10 57 12
rect 11 8 57 10
<< ndif >>
rect 9 24 17 26
rect 9 22 11 24
rect 13 22 17 24
rect 9 20 17 22
rect 19 20 29 26
rect 31 24 39 26
rect 31 22 34 24
rect 36 22 39 24
rect 31 20 39 22
rect 41 24 49 26
rect 41 22 44 24
rect 46 22 49 24
rect 41 20 49 22
rect 51 24 58 26
rect 51 22 54 24
rect 56 22 58 24
rect 51 20 58 22
rect 21 16 27 20
rect 21 14 23 16
rect 25 14 27 16
rect 21 12 27 14
<< pdif >>
rect 53 67 60 69
rect 53 65 55 67
rect 57 65 60 67
rect 37 59 42 65
rect 15 57 22 59
rect 15 55 17 57
rect 19 55 22 57
rect 4 49 9 55
rect 2 47 9 49
rect 2 45 4 47
rect 6 45 9 47
rect 2 43 9 45
rect 11 47 22 55
rect 24 51 32 59
rect 24 49 27 51
rect 29 49 32 51
rect 24 47 32 49
rect 34 57 42 59
rect 34 55 37 57
rect 39 55 42 57
rect 34 47 42 55
rect 44 47 49 65
rect 51 47 60 65
rect 11 43 20 47
<< alu1 >>
rect -2 67 66 72
rect -2 65 5 67
rect 7 65 55 67
rect 57 65 66 67
rect -2 64 66 65
rect 35 57 62 58
rect 35 55 37 57
rect 39 55 62 57
rect 35 54 62 55
rect 17 43 23 50
rect 10 38 23 43
rect 10 36 11 38
rect 13 36 14 38
rect 10 34 14 36
rect 18 33 31 34
rect 18 31 27 33
rect 29 31 31 33
rect 18 30 31 31
rect 18 21 22 30
rect 58 34 62 54
rect 42 30 62 34
rect 42 24 47 30
rect 42 22 44 24
rect 46 22 47 24
rect 42 20 47 22
rect -2 7 66 8
rect -2 5 5 7
rect 7 5 66 7
rect -2 0 66 5
<< ptie >>
rect 3 7 9 9
rect 3 5 5 7
rect 7 5 9 7
rect 3 3 9 5
<< ntie >>
rect 3 67 9 69
rect 3 65 5 67
rect 7 65 9 67
rect 3 63 9 65
<< nmos >>
rect 17 20 19 26
rect 29 20 31 26
rect 39 20 41 26
rect 49 20 51 26
<< pmos >>
rect 9 43 11 55
rect 22 47 24 59
rect 32 47 34 59
rect 42 47 44 65
rect 49 47 51 65
<< polyct0 >>
rect 50 40 52 42
rect 9 14 11 16
rect 57 14 59 16
<< polyct1 >>
rect 11 36 13 38
rect 27 31 29 33
<< ndifct0 >>
rect 11 22 13 24
rect 34 22 36 24
rect 54 22 56 24
rect 23 14 25 16
<< ndifct1 >>
rect 44 22 46 24
<< ntiect1 >>
rect 5 65 7 67
<< ptiect1 >>
rect 5 5 7 7
<< pdifct0 >>
rect 17 55 19 57
rect 4 45 6 47
rect 27 49 29 51
<< pdifct1 >>
rect 55 65 57 67
rect 37 55 39 57
<< alu0 >>
rect 15 57 21 64
rect 15 55 17 57
rect 19 55 21 57
rect 15 54 21 55
rect 26 51 30 53
rect 2 47 7 49
rect 2 45 4 47
rect 6 45 7 47
rect 2 43 7 45
rect 26 49 27 51
rect 29 50 30 51
rect 29 49 38 50
rect 26 46 38 49
rect 2 26 6 43
rect 34 43 38 46
rect 34 42 54 43
rect 34 40 50 42
rect 52 40 54 42
rect 34 39 54 40
rect 2 24 14 26
rect 2 22 11 24
rect 13 22 14 24
rect 7 20 14 22
rect 34 26 38 39
rect 33 24 38 26
rect 33 22 34 24
rect 36 22 38 24
rect 33 20 38 22
rect 53 24 57 26
rect 53 22 54 24
rect 56 22 57 24
rect 7 16 13 20
rect 53 17 57 22
rect 7 14 9 16
rect 11 14 13 16
rect 7 13 13 14
rect 21 16 27 17
rect 21 14 23 16
rect 25 14 27 16
rect 21 8 27 14
rect 53 16 61 17
rect 53 14 57 16
rect 59 14 61 16
rect 53 13 61 14
<< labels >>
rlabel alu0 10 19 10 19 6 bn
rlabel alu0 4 46 4 46 6 bn
rlabel alu0 36 35 36 35 6 an
rlabel alu0 32 48 32 48 6 an
rlabel alu0 55 19 55 19 6 bn
rlabel alu0 44 41 44 41 6 an
rlabel alu1 12 40 12 40 6 b
rlabel polyct1 28 32 28 32 6 a
rlabel alu1 20 24 20 24 6 a
rlabel alu1 20 44 20 44 6 b
rlabel alu1 32 4 32 4 6 vss
rlabel alu1 44 24 44 24 6 z
rlabel alu1 44 56 44 56 6 z
rlabel alu1 32 68 32 68 6 vdd
rlabel alu1 52 32 52 32 6 z
rlabel alu1 60 44 60 44 6 z
rlabel alu1 52 56 52 56 6 z
<< end >>
