magic
tech scmos
timestamp 1552319301
<< nwell >>
rect -5 14 15 30
<< polysilicon >>
rect 2 24 4 26
rect 2 10 4 15
rect 2 3 4 6
rect 2 -5 4 0
<< ndiffusion >>
rect -1 0 2 3
rect 4 0 7 3
<< pdiffusion >>
rect -1 15 2 24
rect 4 15 7 24
<< metal1 >>
rect -5 26 11 30
rect -5 20 -1 26
rect 7 3 11 16
rect -5 -5 -1 -1
rect -5 -9 11 -5
<< ntransistor >>
rect 2 0 4 3
<< ptransistor >>
rect 2 15 4 24
<< polycontact >>
rect 0 6 4 10
<< ndcontact >>
rect -5 -1 -1 3
rect 7 -1 11 3
<< pdcontact >>
rect -5 16 -1 20
rect 7 16 11 20
<< psubstratepcontact >>
rect -9 -9 -5 -5
<< nsubstratencontact >>
rect 11 26 15 30
<< labels >>
rlabel polycontact 2 8 2 8 1 in
rlabel metal1 9 8 9 8 1 out
rlabel metal1 3 28 3 28 5 vdd
rlabel metal1 3 -7 3 -7 1 gnd
<< end >>
