magic
tech scmos
timestamp 1520961445
<< nwell >>
rect -55 -6 13 35
<< polysilicon >>
rect -49 21 -46 23
rect -22 21 -19 23
rect 1 11 4 16
rect -49 -7 -46 5
rect -22 -7 -19 5
rect 1 -7 4 5
rect -47 -11 -46 -7
rect -20 -11 -19 -7
rect 3 -11 4 -7
rect -49 -22 -46 -11
rect -22 -22 -19 -11
rect 1 -22 4 -11
rect -49 -30 -46 -25
rect -22 -30 -19 -25
rect 1 -30 4 -25
<< ndiffusion >>
rect -50 -25 -49 -22
rect -46 -25 -37 -22
rect -33 -25 -22 -22
rect -19 -25 -17 -22
rect -3 -25 1 -22
rect 4 -25 10 -22
<< pdiffusion >>
rect -52 14 -49 21
rect -50 10 -49 14
rect -52 5 -49 10
rect -46 5 -22 21
rect -19 14 -16 21
rect -19 10 -18 14
rect -19 5 -16 10
rect -6 9 1 11
rect -3 5 1 9
rect 4 9 13 11
rect 4 5 9 9
<< metal1 >>
rect -55 27 13 29
rect -55 26 -12 27
rect -54 14 -51 26
rect -8 26 13 27
rect -14 10 -13 13
rect -16 -8 -13 10
rect -5 9 -2 26
rect -3 6 -2 9
rect -16 -11 -1 -8
rect -16 -14 -13 -11
rect -54 -17 -13 -14
rect -54 -21 -51 -17
rect -16 -21 -13 -17
rect 10 -21 13 5
rect -37 -33 -34 -25
rect -7 -33 -4 -25
rect -55 -36 13 -33
<< ntransistor >>
rect -49 -25 -46 -22
rect -22 -25 -19 -22
rect 1 -25 4 -22
<< ptransistor >>
rect -49 5 -46 21
rect -22 5 -19 21
rect 1 5 4 11
<< polycontact >>
rect -51 -11 -47 -7
rect -24 -11 -20 -7
rect -1 -11 3 -7
<< ndcontact >>
rect -54 -25 -50 -21
rect -37 -25 -33 -21
rect -17 -25 -13 -21
rect -7 -25 -3 -21
rect 10 -25 14 -21
<< pdcontact >>
rect -54 10 -50 14
rect -18 10 -14 14
rect -7 5 -3 9
rect 9 5 13 9
<< nsubstratencontact >>
rect -12 23 -8 27
<< labels >>
rlabel metal1 -25 27 -25 27 1 vdd
rlabel polycontact -49 -9 -49 -9 1 A
rlabel polycontact -22 -10 -22 -10 1 B
rlabel pdiffusion -35 12 -35 12 1 n1
rlabel metal1 -36 -35 -36 -35 1 gnd
rlabel metal1 -13 -10 -13 -10 1 or_out
rlabel metal1 11 -10 11 -10 7 out
<< end >>
