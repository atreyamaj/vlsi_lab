* nmos charecteristics varying width working
* with results written to output.txt
*

* device details like model etc.
* include the model files
.include ./t14y_tsmc_025_level3.txt

* spice netlist
m1 drain gate 0 0 cmosn l=3u w=10u


* excitation sources (supply voltages, stimulus etc)
vdd drain 0 dc 5
vgg gate 0 dc 5


* desired responses
.dc vdd 0 5 0.1 vgg 0 5 1


* computing the response for various widths
.control
foreach wid 1.6e-6 6.4e-6 96e-6
* can use any one of the 2 lines below. Both of them give the same result
*alter @m1[w] = $wid
alter m1 w = $wid
run
end
.endc

* plotting the output for various widths
.control
foreach iter 1 2 3  
setplot dc$iter
plot -vdd#branch
end 
.endc

.control
set filetype=ascii
write output.txt 
.endc
.end
