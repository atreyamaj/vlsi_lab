* SPICE3 file created from inverter.ext - technology: scmos

.include ./t14y_tsmc_025_level3.txt

.option scale=1u

M1000 out in vdd vdd cmosp w=6 l=2
+  ad=34 pd=26 as=34 ps=26
M1001 out in gnd Gnd cmosn w=3 l=2
+  ad=25 pd=22 as=25 ps=22
C0 gnd Gnd 3.76fF
C1 in Gnd 4.92fF
Cl out measure 1pF

vsource vdd gnd dc 3.3
vin in gnd dc 3.3 pulse(0 3.3 0 0.1n 0.1n 0.5m 1m)
vcap measure gnd dc 0


.control
dc vin 0 3.3 0.001

meas dc voh find out when in=0.002
meas dc vol find out when in=3.29
let slope=deriv(out)

meas dc vih find in when slope=-1 cross=2
meas dc vil find in when slope=-1 cross=1

let v90 = voh-0.1*(voh-vol)
let v10 = vol+0.1*(voh-vol)
let vhalf = voh-0.5*(voh-vol)

tran 0.1m 4m
plot in out
plot 3.3*vcap#branch
meas tran trise trig out val=dc.v10 rise=1 targ out val=dc.v90 rise=1
meas tran tfall trig out val=dc.v90 fall=1 targ out val=dc.v10 fall=1

meas tran tlh trig in val=1.65 fall=1 targ out val=dc.vhalf rise=1
meas tran thl trig in val=1.65 rise=1 targ out val=dc.vhalf fall=1
let td = 0.5*(thl+tlh)

let power = -3.3*vsource#branch
meas tran pavg AVG power from=0m to=2m 
let pcap = 3.3*abs(vcap#branch)
meas tran pdyn AVG pcap from=0m to=2m

setplot dc1
plot dc1.out
plot deriv(dc1.out)

.endc
.end