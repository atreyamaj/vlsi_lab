* Inverter using a PMOS Transistor varying driver width

.include ./t14y_tsmc_025_level3.txt

* NET List
* m0 drain gate source bulk
m0 out in 0 0 cmosn l=0.25u w=10u
m1 out in supply supply cmosp l=0.25u w=31u
cl out measure 5n

* source
vdd supply 0 dc 3.3
vin in 0 dc 3.3 pulse(0 3.3 0 0.1n 0.1n 0.5m 1m)
vcap measure 0 dc 0


.control
foreach wi 10u 50u
alter @m0[w] = $wi

dc vin 0 3.3 0.001

meas dc voh find out when in=0.002
meas dc vol find out when in=3.29
let slope=deriv(out)

meas dc vih find in when slope=-1 cross=2
meas dc vil find in when slope=-1 cross=1

let v90 = voh-0.1*(voh-vol)
let v10 = vol+0.1*(voh-vol)
let vhalf = voh-0.5*(voh-vol)

tran 0.1m 4m
plot in out
meas tran trise trig out val=dc.v10 rise=1 targ out val=dc.v90 rise=1
meas tran tfall trig out val=dc.v90 fall=1 targ out val=dc.v10 fall=1

meas tran tlh trig in val=1.65 fall=1 targ out val=dc.vhalf rise=1
meas tran thl trig in val=1.65 rise=1 targ out val=dc.vhalf fall=1
let td = 0.5*(thl+tlh)

let power = -3.3*vdd#branch
meas tran pavg AVG power from=0m to=2m 
let pcap = 3.3*abs(vcap#branch)
meas tran pdyn AVG pcap from=0m to=2m
end

setplot dc1
plot dc1.out dc2.out
plot deriv(dc1.out) deriv(dc2.out)
.endc

.end
