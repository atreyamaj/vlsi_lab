* to study NAND gate

.include /home/vlsilab/UG_students_2018/t14y_tsmc_025_level3.txt

Mp1 out ina vdd vdd cmosp l=1u w=2.5u
Mp2 out inb vdd vdd cmosp l=1u w=2.5u
Mn1 out ina n 0 cmosn l=1u w=1u
Mn2 n inb 0 0 cmosn l=1u w=1u

v_dd vdd 0 5
v_a ina 0 PULSE(0 5 0s 0.01ns 0.01ns 3ns 6ns)

v_b inb 0 PULSE(0 5 0s 0.01ns 0.01ns 2.5ns 5ns)



*Trnsfer
.control
*foreach wid 0.1u 1u 10u 100u
*alter Mp1 w = $wid
*alter Mp2 w = $wid
tran 0.01ns 20ns
run

*end
*dc v_a 0 5 0.1

*run
*plot dc1.out deriv(dc1.out) dc2.out deriv(dc2.out) dc3.out deriv(dc3.out) dc4.out deriv(dc4.out)
*plot tran1.out tran2.out tran3.out tran4.out
*meas tran yavg AVG i(v_dd) from=0ns to from= 
plot (out) (vdd*(-v_dd#branch))
*plot 
.endc
.end