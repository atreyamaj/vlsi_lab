magic
tech scmos
timestamp 1552322522
<< nwell >>
rect -5 21 27 23
rect -6 11 27 21
<< polysilicon >>
rect 2 16 4 18
rect 10 16 12 18
rect 2 10 4 13
rect 3 6 4 10
rect 2 3 4 6
rect 10 10 12 13
rect 10 7 21 10
rect 10 3 12 7
rect 2 -2 4 0
rect 10 -2 12 0
<< ndiffusion >>
rect -1 0 2 3
rect 4 0 10 3
rect 12 0 15 3
<< pdiffusion >>
rect -1 13 2 16
rect 4 13 5 16
rect 9 13 10 16
rect 12 13 15 16
<< metal1 >>
rect -5 20 23 23
rect -5 17 -1 20
rect 15 19 23 20
rect 15 17 19 19
rect 6 10 9 13
rect 6 7 18 10
rect 15 3 18 7
rect -5 -4 -1 -1
rect -5 -7 19 -4
<< ntransistor >>
rect 2 0 4 3
rect 10 0 12 3
<< ptransistor >>
rect 2 13 4 16
rect 10 13 12 16
<< polycontact >>
rect -1 6 3 10
rect 21 6 25 10
<< ndcontact >>
rect -5 -1 -1 3
rect 15 -1 19 3
<< pdcontact >>
rect -5 13 -1 17
rect 5 13 9 17
rect 15 13 19 17
<< nsubstratencontact >>
rect 23 19 27 23
<< labels >>
rlabel polycontact 23 8 23 8 7 InA
rlabel polycontact 1 8 1 8 1 InB
rlabel metal1 8 21 8 21 5 Vdd
rlabel metal1 7 -6 7 -6 1 Gnd
rlabel metal1 7 8 7 8 1 Out
<< end >>
