magic
tech scmos
timestamp 1553777430
<< ab >>
rect 0 53 96 67
rect 0 49 2 53
rect 4 49 96 53
rect 0 -5 96 49
<< nwell >>
rect -5 27 101 72
<< pwell >>
rect -5 -10 101 27
<< poly >>
rect 9 61 11 65
rect 32 58 34 63
rect 39 58 41 63
rect 57 61 59 65
rect 67 61 69 65
rect 77 61 79 65
rect 22 49 24 54
rect 9 23 11 36
rect 22 33 24 36
rect 15 31 24 33
rect 15 29 17 31
rect 19 29 21 31
rect 32 30 34 33
rect 39 30 41 33
rect 57 30 59 33
rect 67 30 69 33
rect 77 30 79 33
rect 15 27 21 29
rect 9 21 15 23
rect 9 19 11 21
rect 13 19 15 21
rect 9 17 15 19
rect 9 14 11 17
rect 19 14 21 27
rect 29 28 35 30
rect 29 26 31 28
rect 33 26 35 28
rect 29 24 35 26
rect 39 28 61 30
rect 39 26 50 28
rect 52 26 57 28
rect 59 26 61 28
rect 39 24 61 26
rect 65 28 71 30
rect 65 26 67 28
rect 69 26 71 28
rect 65 24 71 26
rect 75 28 81 30
rect 75 26 77 28
rect 79 26 81 28
rect 75 24 81 26
rect 29 21 31 24
rect 39 21 41 24
rect 59 21 61 24
rect 66 21 68 24
rect 9 -3 11 1
rect 19 -1 21 4
rect 29 2 31 7
rect 39 2 41 7
rect 77 15 79 24
rect 59 -3 61 1
rect 66 -3 68 1
rect 77 -3 79 1
<< ndif >>
rect 24 14 29 21
rect 2 12 9 14
rect 2 10 4 12
rect 6 10 9 12
rect 2 8 9 10
rect 4 1 9 8
rect 11 8 19 14
rect 11 6 14 8
rect 16 6 19 8
rect 11 4 19 6
rect 21 11 29 14
rect 21 9 24 11
rect 26 9 29 11
rect 21 7 29 9
rect 31 19 39 21
rect 31 17 34 19
rect 36 17 39 19
rect 31 7 39 17
rect 41 19 48 21
rect 41 17 44 19
rect 46 17 48 19
rect 41 12 48 17
rect 54 14 59 21
rect 41 10 44 12
rect 46 10 48 12
rect 41 7 48 10
rect 52 12 59 14
rect 52 10 54 12
rect 56 10 59 12
rect 52 8 59 10
rect 21 4 26 7
rect 11 1 16 4
rect 54 1 59 8
rect 61 1 66 21
rect 68 15 75 21
rect 68 5 77 15
rect 68 3 71 5
rect 73 3 77 5
rect 68 1 77 3
rect 79 12 86 15
rect 79 10 82 12
rect 84 10 86 12
rect 79 8 86 10
rect 79 1 84 8
<< pdif >>
rect 4 49 9 61
rect 2 47 9 49
rect 2 45 4 47
rect 6 45 9 47
rect 2 40 9 45
rect 2 38 4 40
rect 6 38 9 40
rect 2 36 9 38
rect 11 59 20 61
rect 11 57 15 59
rect 17 57 20 59
rect 43 59 57 61
rect 43 58 50 59
rect 11 49 20 57
rect 27 49 32 58
rect 11 36 22 49
rect 24 40 32 49
rect 24 38 27 40
rect 29 38 32 40
rect 24 36 32 38
rect 27 33 32 36
rect 34 33 39 58
rect 41 57 50 58
rect 52 57 57 59
rect 41 52 57 57
rect 41 50 50 52
rect 52 50 57 52
rect 41 33 57 50
rect 59 51 67 61
rect 59 49 62 51
rect 64 49 67 51
rect 59 44 67 49
rect 59 42 62 44
rect 64 42 67 44
rect 59 33 67 42
rect 69 59 77 61
rect 69 57 72 59
rect 74 57 77 59
rect 69 52 77 57
rect 69 50 72 52
rect 74 50 77 52
rect 69 33 77 50
rect 79 46 84 61
rect 79 44 86 46
rect 79 42 82 44
rect 84 42 86 44
rect 79 37 86 42
rect 79 35 82 37
rect 84 35 86 37
rect 79 33 86 35
<< alu1 >>
rect -2 59 98 67
rect 2 47 7 49
rect 2 45 4 47
rect 6 45 7 47
rect 2 40 7 45
rect 2 38 4 40
rect 6 38 7 40
rect 2 36 7 38
rect 2 14 6 36
rect 33 33 71 37
rect 33 30 38 33
rect 30 28 38 30
rect 30 26 31 28
rect 33 26 38 28
rect 30 24 38 26
rect 48 28 63 29
rect 48 26 50 28
rect 52 26 57 28
rect 59 26 63 28
rect 48 25 63 26
rect 2 12 7 14
rect 50 16 54 25
rect 81 44 87 46
rect 81 42 82 44
rect 84 42 87 44
rect 81 37 87 42
rect 81 35 82 37
rect 84 35 87 37
rect 81 33 87 35
rect 83 13 87 33
rect 2 10 4 12
rect 6 10 7 12
rect 2 8 7 10
rect 81 12 87 13
rect 81 10 82 12
rect 84 10 87 12
rect 81 9 87 10
rect -2 -5 98 3
<< nmos >>
rect 9 1 11 14
rect 19 4 21 14
rect 29 7 31 21
rect 39 7 41 21
rect 59 1 61 21
rect 66 1 68 21
rect 77 1 79 15
<< pmos >>
rect 9 36 11 61
rect 22 36 24 49
rect 32 33 34 58
rect 39 33 41 58
rect 57 33 59 61
rect 67 33 69 61
rect 77 33 79 61
<< polyct0 >>
rect 17 29 19 31
rect 11 19 13 21
rect 67 26 69 28
rect 77 26 79 28
<< polyct1 >>
rect 31 26 33 28
rect 50 26 52 28
rect 57 26 59 28
<< ndifct0 >>
rect 14 6 16 8
rect 24 9 26 11
rect 34 17 36 19
rect 44 17 46 19
rect 44 10 46 12
rect 54 10 56 12
rect 71 3 73 5
<< ndifct1 >>
rect 4 10 6 12
rect 82 10 84 12
<< pdifct0 >>
rect 15 57 17 59
rect 27 38 29 40
rect 50 57 52 59
rect 50 50 52 52
rect 62 49 64 51
rect 62 42 64 44
rect 72 57 74 59
rect 72 50 74 52
<< pdifct1 >>
rect 4 45 6 47
rect 4 38 6 40
rect 82 42 84 44
rect 82 35 84 37
<< alu0 >>
rect 13 57 15 59
rect 17 57 19 59
rect 13 56 19 57
rect 48 57 50 59
rect 52 57 54 59
rect 48 52 54 57
rect 70 57 72 59
rect 74 57 76 59
rect 48 50 50 52
rect 52 50 54 52
rect 48 49 54 50
rect 61 51 65 53
rect 61 49 62 51
rect 64 49 65 51
rect 70 52 76 57
rect 70 50 72 52
rect 74 50 76 52
rect 70 49 76 50
rect 18 45 42 49
rect 61 45 65 49
rect 16 41 22 45
rect 38 44 78 45
rect 38 42 62 44
rect 64 42 78 44
rect 16 31 20 41
rect 26 40 30 42
rect 38 41 78 42
rect 26 38 27 40
rect 29 38 30 40
rect 26 37 30 38
rect 16 29 17 31
rect 19 29 20 31
rect 16 27 20 29
rect 23 33 30 37
rect 23 22 27 33
rect 66 28 70 33
rect 66 26 67 28
rect 69 26 70 28
rect 9 21 27 22
rect 9 19 11 21
rect 13 20 27 21
rect 13 19 38 20
rect 9 18 34 19
rect 23 17 34 18
rect 36 17 38 19
rect 23 16 38 17
rect 43 19 47 21
rect 43 17 44 19
rect 46 17 47 19
rect 43 12 47 17
rect 66 24 70 26
rect 74 30 78 41
rect 74 28 80 30
rect 74 26 77 28
rect 79 26 80 28
rect 74 24 80 26
rect 74 21 78 24
rect 58 17 78 21
rect 58 13 62 17
rect 22 11 44 12
rect 13 8 17 10
rect 22 9 24 11
rect 26 10 44 11
rect 46 10 47 12
rect 26 9 47 10
rect 52 12 62 13
rect 52 10 54 12
rect 56 10 62 12
rect 52 9 62 10
rect 22 8 47 9
rect 13 6 14 8
rect 16 6 17 8
rect 13 3 17 6
rect 69 5 75 6
rect 69 3 71 5
rect 73 3 75 5
<< labels >>
rlabel alu1 4 27 4 27 6 so
rlabel alu1 48 63 48 63 6 vdd
rlabel alu1 84 39 84 39 6 co
rlabel alu1 48 -1 48 -1 1 gnd
rlabel alu1 60 27 60 27 6 a
rlabel alu1 52 35 52 35 1 b
<< end >>
