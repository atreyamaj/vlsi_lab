* SPICE3 file created from aoi.ext - technology: scmos

.include /home/vlsilab/UG_students_2018/t14y_tsmc_025_level3.txt

M1000 vdd B n2 vdd cmosp w=12u l=2u
+  ad=108p pd=42u as=132p ps=74u
M1001 n2 C vdd vdd cmosp w=12u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1002 out A n2 vdd cmosp w=12u l=2u
+  ad=96p pd=40u as=0p ps=0u
M1003 n1 B out Gnd cmosn w=6u l=2u
+  ad=54p pd=30u as=54p ps=46u
M1004 gnd C n1 Gnd cmosn w=6u l=2u
+  ad=39p pd=26u as=0p ps=0u
M1005 out A gnd Gnd cmosn w=3u l=2u
+  ad=0p pd=0u as=0p ps=0u

C0 gnd Gnd 3.29fF
C1 out Gnd 6.58fF
C2 n2 Gnd 3.06fF
C3 A Gnd 6.59fF
C4 C Gnd 6.19fF
C5 B Gnd 6.19fF

v_dd vdd 0 5
gd gnd 0 0 

v_ina A 0 PULSE(0 5 0 0.1n 0.1n 50n 100n)
v_inb B 0 PULSE(0 5 0 0.1n 0.1n 40n 80n)
v_inc C 0 PULSE(0 5 0 0.1n 0.1n 30n 60n)


.control
tran 0.1n 300n
run
plot (out) (0.125*A) (0.25*B) (0.5*C)

.endc

.end
