magic
tech scmos
timestamp 1553798959
<< rotate >>
rect 97 -65 108 -63
rect 74 -69 76 -67
rect 97 -72 111 -65
rect 100 -74 111 -72
<< ab >>
rect 27 58 204 72
rect 27 54 29 58
rect 31 54 201 58
rect 203 54 204 58
rect 27 -54 204 54
rect 27 -58 29 -54
rect 31 -58 201 -54
rect 203 -58 204 -54
rect 27 -72 204 -58
rect 206 -39 247 72
rect 206 -42 248 -39
rect 206 -72 247 -42
<< nwell >>
rect 22 32 250 77
rect 22 -77 250 -32
<< pwell >>
rect 22 -32 250 32
<< poly >>
rect 36 66 38 70
rect 59 63 61 68
rect 66 63 68 68
rect 84 66 86 70
rect 94 66 96 70
rect 104 66 106 70
rect 126 66 128 70
rect 136 66 138 70
rect 146 66 148 70
rect 49 54 51 59
rect 36 28 38 41
rect 49 38 51 41
rect 164 63 166 68
rect 171 63 173 68
rect 194 66 196 70
rect 215 66 217 70
rect 222 66 224 70
rect 181 54 183 59
rect 235 56 237 61
rect 215 42 217 45
rect 181 38 183 41
rect 42 36 51 38
rect 42 34 44 36
rect 46 34 48 36
rect 59 35 61 38
rect 66 35 68 38
rect 84 35 86 38
rect 94 35 96 38
rect 104 35 106 38
rect 126 35 128 38
rect 136 35 138 38
rect 146 35 148 38
rect 164 35 166 38
rect 171 35 173 38
rect 181 36 190 38
rect 42 32 48 34
rect 36 26 42 28
rect 36 24 38 26
rect 40 24 42 26
rect 36 22 42 24
rect 36 19 38 22
rect 46 19 48 32
rect 56 33 62 35
rect 56 31 58 33
rect 60 31 62 33
rect 56 29 62 31
rect 66 33 88 35
rect 66 31 77 33
rect 79 31 84 33
rect 86 31 88 33
rect 66 29 88 31
rect 92 33 98 35
rect 92 31 94 33
rect 96 31 98 33
rect 92 29 98 31
rect 102 33 108 35
rect 102 31 104 33
rect 106 31 108 33
rect 102 29 108 31
rect 124 33 130 35
rect 124 31 126 33
rect 128 31 130 33
rect 124 29 130 31
rect 134 33 140 35
rect 134 31 136 33
rect 138 31 140 33
rect 134 29 140 31
rect 144 33 166 35
rect 144 31 146 33
rect 148 31 153 33
rect 155 31 166 33
rect 144 29 166 31
rect 170 33 176 35
rect 170 31 172 33
rect 174 31 176 33
rect 170 29 176 31
rect 56 26 58 29
rect 66 26 68 29
rect 86 26 88 29
rect 93 26 95 29
rect 36 2 38 6
rect 46 4 48 9
rect 56 7 58 12
rect 66 7 68 12
rect 104 20 106 29
rect 126 20 128 29
rect 137 26 139 29
rect 144 26 146 29
rect 164 26 166 29
rect 174 26 176 29
rect 184 34 186 36
rect 188 34 190 36
rect 184 32 190 34
rect 184 19 186 32
rect 194 28 196 41
rect 211 40 217 42
rect 211 38 213 40
rect 215 38 217 40
rect 211 36 217 38
rect 190 26 196 28
rect 215 26 217 36
rect 222 35 224 45
rect 235 35 237 38
rect 221 33 227 35
rect 221 31 223 33
rect 225 31 227 33
rect 221 29 227 31
rect 231 33 237 35
rect 231 31 233 33
rect 235 31 237 33
rect 231 29 237 31
rect 225 26 227 29
rect 235 26 237 29
rect 190 24 192 26
rect 194 24 196 26
rect 190 22 196 24
rect 194 19 196 22
rect 164 7 166 12
rect 174 7 176 12
rect 86 2 88 6
rect 93 2 95 6
rect 104 2 106 6
rect 126 2 128 6
rect 137 2 139 6
rect 144 2 146 6
rect 184 4 186 9
rect 215 15 217 20
rect 225 15 227 20
rect 235 12 237 17
rect 194 2 196 6
rect 36 -6 38 -2
rect 46 -9 48 -4
rect 86 -6 88 -2
rect 93 -6 95 -2
rect 104 -6 106 -2
rect 126 -6 128 -2
rect 137 -6 139 -2
rect 144 -6 146 -2
rect 56 -12 58 -7
rect 66 -12 68 -7
rect 36 -22 38 -19
rect 36 -24 42 -22
rect 36 -26 38 -24
rect 40 -26 42 -24
rect 36 -28 42 -26
rect 36 -41 38 -28
rect 46 -32 48 -19
rect 42 -34 48 -32
rect 42 -36 44 -34
rect 46 -36 48 -34
rect 56 -29 58 -26
rect 66 -29 68 -26
rect 86 -29 88 -26
rect 93 -29 95 -26
rect 104 -29 106 -20
rect 126 -29 128 -20
rect 164 -12 166 -7
rect 174 -12 176 -7
rect 184 -9 186 -4
rect 194 -6 196 -2
rect 137 -29 139 -26
rect 144 -29 146 -26
rect 164 -29 166 -26
rect 174 -29 176 -26
rect 56 -31 62 -29
rect 56 -33 58 -31
rect 60 -33 62 -31
rect 56 -35 62 -33
rect 66 -31 88 -29
rect 66 -33 77 -31
rect 79 -33 84 -31
rect 86 -33 88 -31
rect 66 -35 88 -33
rect 92 -31 98 -29
rect 92 -33 94 -31
rect 96 -33 98 -31
rect 92 -35 98 -33
rect 102 -31 108 -29
rect 102 -33 104 -31
rect 106 -33 108 -31
rect 102 -35 108 -33
rect 124 -31 130 -29
rect 124 -33 126 -31
rect 128 -33 130 -31
rect 124 -35 130 -33
rect 134 -31 140 -29
rect 134 -33 136 -31
rect 138 -33 140 -31
rect 134 -35 140 -33
rect 144 -31 166 -29
rect 144 -33 146 -31
rect 148 -33 153 -31
rect 155 -33 166 -31
rect 144 -35 166 -33
rect 170 -31 176 -29
rect 170 -33 172 -31
rect 174 -33 176 -31
rect 170 -35 176 -33
rect 184 -32 186 -19
rect 194 -22 196 -19
rect 190 -24 196 -22
rect 190 -26 192 -24
rect 194 -26 196 -24
rect 215 -20 217 -15
rect 225 -20 227 -15
rect 235 -17 237 -12
rect 190 -28 196 -26
rect 184 -34 190 -32
rect 42 -38 51 -36
rect 59 -38 61 -35
rect 66 -38 68 -35
rect 84 -38 86 -35
rect 94 -38 96 -35
rect 104 -38 106 -35
rect 126 -38 128 -35
rect 136 -38 138 -35
rect 146 -38 148 -35
rect 164 -38 166 -35
rect 171 -38 173 -35
rect 184 -36 186 -34
rect 188 -36 190 -34
rect 181 -38 190 -36
rect 49 -41 51 -38
rect 49 -59 51 -54
rect 36 -70 38 -66
rect 59 -68 61 -63
rect 66 -68 68 -63
rect 181 -41 183 -38
rect 194 -41 196 -28
rect 215 -36 217 -26
rect 225 -29 227 -26
rect 235 -29 237 -26
rect 221 -31 227 -29
rect 221 -33 223 -31
rect 225 -33 227 -31
rect 221 -35 227 -33
rect 231 -31 237 -29
rect 231 -33 233 -31
rect 235 -33 237 -31
rect 231 -35 237 -33
rect 211 -38 217 -36
rect 211 -40 213 -38
rect 215 -40 217 -38
rect 181 -59 183 -54
rect 84 -70 86 -66
rect 94 -70 96 -66
rect 104 -70 106 -66
rect 126 -70 128 -66
rect 136 -70 138 -66
rect 146 -70 148 -66
rect 164 -68 166 -63
rect 171 -68 173 -63
rect 211 -42 217 -40
rect 215 -45 217 -42
rect 222 -45 224 -35
rect 235 -38 237 -35
rect 235 -61 237 -56
rect 194 -70 196 -66
rect 215 -70 217 -66
rect 222 -70 224 -66
<< ndif >>
rect 51 19 56 26
rect 29 17 36 19
rect 29 15 31 17
rect 33 15 36 17
rect 29 13 36 15
rect 31 6 36 13
rect 38 13 46 19
rect 38 11 41 13
rect 43 11 46 13
rect 38 9 46 11
rect 48 16 56 19
rect 48 14 51 16
rect 53 14 56 16
rect 48 12 56 14
rect 58 24 66 26
rect 58 22 61 24
rect 63 22 66 24
rect 58 12 66 22
rect 68 24 75 26
rect 68 22 71 24
rect 73 22 75 24
rect 68 17 75 22
rect 81 19 86 26
rect 68 15 71 17
rect 73 15 75 17
rect 68 12 75 15
rect 79 17 86 19
rect 79 15 81 17
rect 83 15 86 17
rect 79 13 86 15
rect 48 9 53 12
rect 38 6 43 9
rect 81 6 86 13
rect 88 6 93 26
rect 95 20 102 26
rect 130 20 137 26
rect 95 10 104 20
rect 95 8 98 10
rect 100 8 104 10
rect 95 6 104 8
rect 106 17 113 20
rect 106 15 109 17
rect 111 15 113 17
rect 106 13 113 15
rect 119 17 126 20
rect 119 15 121 17
rect 123 15 126 17
rect 119 13 126 15
rect 106 6 111 13
rect 121 6 126 13
rect 128 10 137 20
rect 128 8 132 10
rect 134 8 137 10
rect 128 6 137 8
rect 139 6 144 26
rect 146 19 151 26
rect 157 24 164 26
rect 157 22 159 24
rect 161 22 164 24
rect 146 17 153 19
rect 146 15 149 17
rect 151 15 153 17
rect 146 13 153 15
rect 157 17 164 22
rect 157 15 159 17
rect 161 15 164 17
rect 146 6 151 13
rect 157 12 164 15
rect 166 24 174 26
rect 166 22 169 24
rect 171 22 174 24
rect 166 12 174 22
rect 176 19 181 26
rect 208 20 215 26
rect 217 24 225 26
rect 217 22 220 24
rect 222 22 225 24
rect 217 20 225 22
rect 227 20 235 26
rect 176 16 184 19
rect 176 14 179 16
rect 181 14 184 16
rect 176 12 184 14
rect 179 9 184 12
rect 186 13 194 19
rect 186 11 189 13
rect 191 11 194 13
rect 186 9 194 11
rect 189 6 194 9
rect 196 17 203 19
rect 196 15 199 17
rect 201 15 203 17
rect 196 13 203 15
rect 208 13 213 20
rect 229 17 235 20
rect 237 24 244 26
rect 237 22 240 24
rect 242 22 244 24
rect 237 20 244 22
rect 237 17 242 20
rect 229 13 233 17
rect 196 6 201 13
rect 208 11 214 13
rect 208 9 210 11
rect 212 9 214 11
rect 208 7 214 9
rect 227 11 233 13
rect 227 9 229 11
rect 231 9 233 11
rect 227 7 233 9
rect 31 -13 36 -6
rect 29 -15 36 -13
rect 29 -17 31 -15
rect 33 -17 36 -15
rect 29 -19 36 -17
rect 38 -9 43 -6
rect 38 -11 46 -9
rect 38 -13 41 -11
rect 43 -13 46 -11
rect 38 -19 46 -13
rect 48 -12 53 -9
rect 48 -14 56 -12
rect 48 -16 51 -14
rect 53 -16 56 -14
rect 48 -19 56 -16
rect 51 -26 56 -19
rect 58 -22 66 -12
rect 58 -24 61 -22
rect 63 -24 66 -22
rect 58 -26 66 -24
rect 68 -15 75 -12
rect 81 -13 86 -6
rect 68 -17 71 -15
rect 73 -17 75 -15
rect 68 -22 75 -17
rect 79 -15 86 -13
rect 79 -17 81 -15
rect 83 -17 86 -15
rect 79 -19 86 -17
rect 68 -24 71 -22
rect 73 -24 75 -22
rect 68 -26 75 -24
rect 81 -26 86 -19
rect 88 -26 93 -6
rect 95 -8 104 -6
rect 95 -10 98 -8
rect 100 -10 104 -8
rect 95 -20 104 -10
rect 106 -13 111 -6
rect 121 -13 126 -6
rect 106 -15 113 -13
rect 106 -17 109 -15
rect 111 -17 113 -15
rect 106 -20 113 -17
rect 119 -15 126 -13
rect 119 -17 121 -15
rect 123 -17 126 -15
rect 119 -20 126 -17
rect 128 -8 137 -6
rect 128 -10 132 -8
rect 134 -10 137 -8
rect 128 -20 137 -10
rect 95 -26 102 -20
rect 130 -26 137 -20
rect 139 -26 144 -6
rect 146 -13 151 -6
rect 189 -9 194 -6
rect 179 -12 184 -9
rect 146 -15 153 -13
rect 146 -17 149 -15
rect 151 -17 153 -15
rect 146 -19 153 -17
rect 157 -15 164 -12
rect 157 -17 159 -15
rect 161 -17 164 -15
rect 146 -26 151 -19
rect 157 -22 164 -17
rect 157 -24 159 -22
rect 161 -24 164 -22
rect 157 -26 164 -24
rect 166 -22 174 -12
rect 166 -24 169 -22
rect 171 -24 174 -22
rect 166 -26 174 -24
rect 176 -14 184 -12
rect 176 -16 179 -14
rect 181 -16 184 -14
rect 176 -19 184 -16
rect 186 -11 194 -9
rect 186 -13 189 -11
rect 191 -13 194 -11
rect 186 -19 194 -13
rect 196 -13 201 -6
rect 208 -9 214 -7
rect 208 -11 210 -9
rect 212 -11 214 -9
rect 208 -13 214 -11
rect 227 -9 233 -7
rect 227 -11 229 -9
rect 231 -11 233 -9
rect 227 -13 233 -11
rect 196 -15 203 -13
rect 196 -17 199 -15
rect 201 -17 203 -15
rect 196 -19 203 -17
rect 176 -26 181 -19
rect 208 -20 213 -13
rect 229 -17 233 -13
rect 229 -20 235 -17
rect 208 -26 215 -20
rect 217 -22 225 -20
rect 217 -24 220 -22
rect 222 -24 225 -22
rect 217 -26 225 -24
rect 227 -26 235 -20
rect 237 -20 242 -17
rect 237 -22 244 -20
rect 237 -24 240 -22
rect 242 -24 244 -22
rect 237 -26 244 -24
<< pdif >>
rect 31 54 36 66
rect 29 52 36 54
rect 29 50 31 52
rect 33 50 36 52
rect 29 45 36 50
rect 29 43 31 45
rect 33 43 36 45
rect 29 41 36 43
rect 38 64 47 66
rect 38 62 42 64
rect 44 62 47 64
rect 70 64 84 66
rect 70 63 77 64
rect 38 54 47 62
rect 54 54 59 63
rect 38 41 49 54
rect 51 45 59 54
rect 51 43 54 45
rect 56 43 59 45
rect 51 41 59 43
rect 54 38 59 41
rect 61 38 66 63
rect 68 62 77 63
rect 79 62 84 64
rect 68 57 84 62
rect 68 55 77 57
rect 79 55 84 57
rect 68 38 84 55
rect 86 56 94 66
rect 86 54 89 56
rect 91 54 94 56
rect 86 49 94 54
rect 86 47 89 49
rect 91 47 94 49
rect 86 38 94 47
rect 96 64 104 66
rect 96 62 99 64
rect 101 62 104 64
rect 96 57 104 62
rect 96 55 99 57
rect 101 55 104 57
rect 96 38 104 55
rect 106 51 111 66
rect 121 51 126 66
rect 106 49 113 51
rect 106 47 109 49
rect 111 47 113 49
rect 106 42 113 47
rect 106 40 109 42
rect 111 40 113 42
rect 106 38 113 40
rect 119 49 126 51
rect 119 47 121 49
rect 123 47 126 49
rect 119 42 126 47
rect 119 40 121 42
rect 123 40 126 42
rect 119 38 126 40
rect 128 64 136 66
rect 128 62 131 64
rect 133 62 136 64
rect 128 57 136 62
rect 128 55 131 57
rect 133 55 136 57
rect 128 38 136 55
rect 138 56 146 66
rect 138 54 141 56
rect 143 54 146 56
rect 138 49 146 54
rect 138 47 141 49
rect 143 47 146 49
rect 138 38 146 47
rect 148 64 162 66
rect 148 62 153 64
rect 155 63 162 64
rect 185 64 194 66
rect 155 62 164 63
rect 148 57 164 62
rect 148 55 153 57
rect 155 55 164 57
rect 148 38 164 55
rect 166 38 171 63
rect 173 54 178 63
rect 185 62 188 64
rect 190 62 194 64
rect 185 54 194 62
rect 173 45 181 54
rect 173 43 176 45
rect 178 43 181 45
rect 173 41 181 43
rect 183 41 194 54
rect 196 54 201 66
rect 210 59 215 66
rect 208 57 215 59
rect 208 55 210 57
rect 212 55 215 57
rect 196 52 203 54
rect 208 53 215 55
rect 196 50 199 52
rect 201 50 203 52
rect 196 45 203 50
rect 210 45 215 53
rect 217 45 222 66
rect 224 64 233 66
rect 224 62 229 64
rect 231 62 233 64
rect 224 56 233 62
rect 224 45 235 56
rect 196 43 199 45
rect 201 43 203 45
rect 196 41 203 43
rect 173 38 178 41
rect 227 38 235 45
rect 237 54 244 56
rect 237 52 240 54
rect 242 52 244 54
rect 237 47 244 52
rect 237 45 240 47
rect 242 45 244 47
rect 237 43 244 45
rect 237 38 242 43
rect 54 -41 59 -38
rect 29 -43 36 -41
rect 29 -45 31 -43
rect 33 -45 36 -43
rect 29 -50 36 -45
rect 29 -52 31 -50
rect 33 -52 36 -50
rect 29 -54 36 -52
rect 31 -66 36 -54
rect 38 -54 49 -41
rect 51 -43 59 -41
rect 51 -45 54 -43
rect 56 -45 59 -43
rect 51 -54 59 -45
rect 38 -62 47 -54
rect 38 -64 42 -62
rect 44 -64 47 -62
rect 54 -63 59 -54
rect 61 -63 66 -38
rect 68 -55 84 -38
rect 68 -57 77 -55
rect 79 -57 84 -55
rect 68 -62 84 -57
rect 68 -63 77 -62
rect 38 -66 47 -64
rect 70 -64 77 -63
rect 79 -64 84 -62
rect 70 -66 84 -64
rect 86 -47 94 -38
rect 86 -49 89 -47
rect 91 -49 94 -47
rect 86 -54 94 -49
rect 86 -56 89 -54
rect 91 -56 94 -54
rect 86 -66 94 -56
rect 96 -55 104 -38
rect 96 -57 99 -55
rect 101 -57 104 -55
rect 96 -62 104 -57
rect 96 -64 99 -62
rect 101 -64 104 -62
rect 96 -66 104 -64
rect 106 -40 113 -38
rect 106 -42 109 -40
rect 111 -42 113 -40
rect 106 -47 113 -42
rect 106 -49 109 -47
rect 111 -49 113 -47
rect 106 -51 113 -49
rect 119 -40 126 -38
rect 119 -42 121 -40
rect 123 -42 126 -40
rect 119 -47 126 -42
rect 119 -49 121 -47
rect 123 -49 126 -47
rect 119 -51 126 -49
rect 106 -66 111 -51
rect 121 -66 126 -51
rect 128 -55 136 -38
rect 128 -57 131 -55
rect 133 -57 136 -55
rect 128 -62 136 -57
rect 128 -64 131 -62
rect 133 -64 136 -62
rect 128 -66 136 -64
rect 138 -47 146 -38
rect 138 -49 141 -47
rect 143 -49 146 -47
rect 138 -54 146 -49
rect 138 -56 141 -54
rect 143 -56 146 -54
rect 138 -66 146 -56
rect 148 -55 164 -38
rect 148 -57 153 -55
rect 155 -57 164 -55
rect 148 -62 164 -57
rect 148 -64 153 -62
rect 155 -63 164 -62
rect 166 -63 171 -38
rect 173 -41 178 -38
rect 173 -43 181 -41
rect 173 -45 176 -43
rect 178 -45 181 -43
rect 173 -54 181 -45
rect 183 -54 194 -41
rect 173 -63 178 -54
rect 185 -62 194 -54
rect 155 -64 162 -63
rect 148 -66 162 -64
rect 185 -64 188 -62
rect 190 -64 194 -62
rect 185 -66 194 -64
rect 196 -43 203 -41
rect 196 -45 199 -43
rect 201 -45 203 -43
rect 227 -45 235 -38
rect 196 -50 203 -45
rect 196 -52 199 -50
rect 201 -52 203 -50
rect 196 -54 203 -52
rect 210 -53 215 -45
rect 196 -66 201 -54
rect 208 -55 215 -53
rect 208 -57 210 -55
rect 212 -57 215 -55
rect 208 -59 215 -57
rect 210 -66 215 -59
rect 217 -66 222 -45
rect 224 -56 235 -45
rect 237 -43 242 -38
rect 237 -45 244 -43
rect 237 -47 240 -45
rect 242 -47 244 -45
rect 237 -52 244 -47
rect 237 -54 240 -52
rect 242 -54 244 -52
rect 237 -56 244 -54
rect 224 -62 233 -56
rect 224 -64 229 -62
rect 231 -64 233 -62
rect 224 -66 233 -64
<< alu1 >>
rect 25 67 247 72
rect 25 65 239 67
rect 241 65 247 67
rect 25 64 247 65
rect 240 58 244 59
rect 231 54 244 58
rect 29 52 34 54
rect 29 50 31 52
rect 33 50 34 52
rect 29 45 34 50
rect 29 43 31 45
rect 33 43 34 45
rect 29 41 34 43
rect 29 25 33 41
rect 60 38 98 42
rect 60 35 65 38
rect 57 33 65 35
rect 57 31 58 33
rect 60 31 65 33
rect 57 29 65 31
rect 75 33 90 34
rect 75 31 77 33
rect 79 31 84 33
rect 86 31 90 33
rect 75 30 90 31
rect 29 23 30 25
rect 32 23 33 25
rect 29 19 33 23
rect 29 17 34 19
rect 77 21 81 30
rect 108 49 114 51
rect 108 47 109 49
rect 111 47 114 49
rect 108 42 114 47
rect 108 40 109 42
rect 111 40 114 42
rect 108 38 114 40
rect 110 33 114 38
rect 110 31 111 33
rect 113 31 114 33
rect 110 18 114 31
rect 29 15 31 17
rect 33 15 34 17
rect 29 13 34 15
rect 108 17 114 18
rect 108 15 109 17
rect 111 15 114 17
rect 108 14 114 15
rect 118 49 124 51
rect 198 52 203 54
rect 198 50 199 52
rect 201 50 203 52
rect 118 47 121 49
rect 123 47 124 49
rect 118 46 124 47
rect 118 44 121 46
rect 123 44 124 46
rect 118 42 124 44
rect 118 40 121 42
rect 123 40 124 42
rect 118 38 124 40
rect 118 18 122 38
rect 134 38 172 42
rect 167 35 172 38
rect 142 33 157 34
rect 142 31 146 33
rect 148 31 153 33
rect 155 31 157 33
rect 142 30 157 31
rect 167 33 175 35
rect 167 31 172 33
rect 174 31 175 33
rect 151 25 155 30
rect 167 29 175 31
rect 198 45 203 50
rect 198 43 199 45
rect 201 43 203 45
rect 198 41 203 43
rect 151 23 152 25
rect 154 23 155 25
rect 151 21 155 23
rect 118 17 124 18
rect 118 15 121 17
rect 123 15 124 17
rect 118 14 124 15
rect 199 19 203 41
rect 208 46 212 51
rect 208 44 209 46
rect 211 44 212 46
rect 208 42 212 44
rect 208 40 229 42
rect 208 38 213 40
rect 215 38 229 40
rect 208 33 229 34
rect 208 31 209 33
rect 211 31 223 33
rect 225 31 229 33
rect 208 30 229 31
rect 242 52 244 54
rect 240 47 244 52
rect 242 45 244 47
rect 208 21 212 30
rect 240 29 244 45
rect 240 27 241 29
rect 243 27 244 29
rect 240 26 244 27
rect 239 24 244 26
rect 239 22 240 24
rect 242 22 244 24
rect 239 20 244 22
rect 198 17 203 19
rect 198 15 199 17
rect 201 15 203 17
rect 198 13 203 15
rect 25 7 247 8
rect 25 5 239 7
rect 241 5 247 7
rect 25 -5 247 5
rect 25 -7 239 -5
rect 241 -7 247 -5
rect 25 -8 247 -7
rect 29 -15 34 -13
rect 29 -17 31 -15
rect 33 -17 34 -15
rect 29 -19 34 -17
rect 29 -23 33 -19
rect 29 -25 30 -23
rect 32 -25 33 -23
rect 29 -41 33 -25
rect 108 -15 114 -14
rect 108 -17 109 -15
rect 111 -17 114 -15
rect 108 -18 114 -17
rect 29 -43 34 -41
rect 29 -45 31 -43
rect 33 -45 34 -43
rect 29 -50 34 -45
rect 57 -31 65 -29
rect 77 -30 81 -21
rect 57 -33 58 -31
rect 60 -33 65 -31
rect 57 -35 65 -33
rect 75 -31 90 -30
rect 75 -33 77 -31
rect 79 -33 84 -31
rect 86 -33 90 -31
rect 75 -34 90 -33
rect 60 -38 65 -35
rect 110 -31 114 -18
rect 110 -33 111 -31
rect 113 -33 114 -31
rect 60 -42 98 -38
rect 110 -38 114 -33
rect 108 -40 114 -38
rect 108 -42 109 -40
rect 111 -42 114 -40
rect 108 -47 114 -42
rect 108 -49 109 -47
rect 111 -49 114 -47
rect 29 -52 31 -50
rect 33 -52 34 -50
rect 29 -54 34 -52
rect 108 -51 114 -49
rect 118 -15 124 -14
rect 118 -17 121 -15
rect 123 -17 124 -15
rect 118 -18 124 -17
rect 198 -15 203 -13
rect 198 -17 199 -15
rect 201 -17 203 -15
rect 118 -38 122 -18
rect 151 -23 155 -21
rect 151 -25 152 -23
rect 154 -25 155 -23
rect 118 -40 124 -38
rect 118 -42 121 -40
rect 123 -42 124 -40
rect 118 -44 124 -42
rect 118 -46 121 -44
rect 123 -46 124 -44
rect 118 -47 124 -46
rect 118 -49 121 -47
rect 123 -49 124 -47
rect 118 -51 124 -49
rect 151 -30 155 -25
rect 198 -19 203 -17
rect 142 -31 157 -30
rect 142 -33 146 -31
rect 148 -33 153 -31
rect 155 -33 157 -31
rect 142 -34 157 -33
rect 167 -31 175 -29
rect 167 -33 172 -31
rect 174 -33 175 -31
rect 167 -35 175 -33
rect 167 -36 172 -35
rect 167 -38 169 -36
rect 171 -38 172 -36
rect 134 -42 172 -38
rect 199 -41 203 -19
rect 208 -25 212 -21
rect 208 -27 209 -25
rect 211 -27 212 -25
rect 208 -30 212 -27
rect 208 -31 229 -30
rect 208 -33 223 -31
rect 225 -33 229 -31
rect 208 -34 229 -33
rect 239 -22 244 -20
rect 239 -24 240 -22
rect 242 -24 244 -22
rect 239 -26 244 -24
rect 198 -43 203 -41
rect 198 -45 199 -43
rect 201 -45 203 -43
rect 198 -50 203 -45
rect 198 -52 199 -50
rect 201 -52 203 -50
rect 208 -40 213 -38
rect 215 -40 229 -38
rect 208 -42 229 -40
rect 208 -44 212 -42
rect 208 -46 209 -44
rect 211 -46 212 -44
rect 208 -51 212 -46
rect 198 -54 203 -52
rect 240 -45 244 -26
rect 242 -47 244 -45
rect 240 -52 244 -47
rect 242 -54 244 -52
rect 231 -58 244 -54
rect 240 -59 244 -58
rect 25 -65 247 -64
rect 25 -67 239 -65
rect 241 -67 247 -65
rect 25 -72 247 -67
<< alu2 >>
rect 120 46 212 47
rect 120 44 121 46
rect 123 44 209 46
rect 211 44 212 46
rect 120 43 212 44
rect 110 33 213 34
rect 110 31 111 33
rect 113 31 209 33
rect 211 31 213 33
rect 110 30 213 31
rect 240 29 248 30
rect 240 27 241 29
rect 243 27 245 29
rect 247 27 248 29
rect 240 26 248 27
rect 29 25 155 26
rect 29 23 30 25
rect 32 23 152 25
rect 154 23 155 25
rect 29 22 155 23
rect 29 -23 155 -22
rect 29 -25 30 -23
rect 32 -25 152 -23
rect 154 -25 155 -23
rect 29 -26 155 -25
rect 159 -25 212 -24
rect 159 -27 209 -25
rect 211 -27 212 -25
rect 159 -28 212 -27
rect 159 -30 163 -28
rect 110 -31 163 -30
rect 110 -33 111 -31
rect 113 -33 163 -31
rect 110 -34 163 -33
rect 168 -36 248 -35
rect 168 -38 169 -36
rect 171 -38 245 -36
rect 247 -38 248 -36
rect 168 -39 248 -38
rect 120 -44 212 -43
rect 120 -46 121 -44
rect 123 -46 209 -44
rect 211 -46 212 -44
rect 120 -47 212 -46
<< alu3 >>
rect 244 29 248 30
rect 244 27 245 29
rect 247 27 248 29
rect 244 -36 248 27
rect 244 -38 245 -36
rect 247 -38 248 -36
rect 244 -39 248 -38
<< ptie >>
rect 237 7 243 9
rect 237 5 239 7
rect 241 5 243 7
rect 237 3 243 5
rect 237 -5 243 -3
rect 237 -7 239 -5
rect 241 -7 243 -5
rect 237 -9 243 -7
<< ntie >>
rect 237 67 243 69
rect 237 65 239 67
rect 241 65 243 67
rect 237 63 243 65
rect 237 -65 243 -63
rect 237 -67 239 -65
rect 241 -67 243 -65
rect 237 -69 243 -67
<< nmos >>
rect 36 6 38 19
rect 46 9 48 19
rect 56 12 58 26
rect 66 12 68 26
rect 86 6 88 26
rect 93 6 95 26
rect 104 6 106 20
rect 126 6 128 20
rect 137 6 139 26
rect 144 6 146 26
rect 164 12 166 26
rect 174 12 176 26
rect 215 20 217 26
rect 225 20 227 26
rect 184 9 186 19
rect 194 6 196 19
rect 235 17 237 26
rect 36 -19 38 -6
rect 46 -19 48 -9
rect 56 -26 58 -12
rect 66 -26 68 -12
rect 86 -26 88 -6
rect 93 -26 95 -6
rect 104 -20 106 -6
rect 126 -20 128 -6
rect 137 -26 139 -6
rect 144 -26 146 -6
rect 164 -26 166 -12
rect 174 -26 176 -12
rect 184 -19 186 -9
rect 194 -19 196 -6
rect 215 -26 217 -20
rect 225 -26 227 -20
rect 235 -26 237 -17
<< pmos >>
rect 36 41 38 66
rect 49 41 51 54
rect 59 38 61 63
rect 66 38 68 63
rect 84 38 86 66
rect 94 38 96 66
rect 104 38 106 66
rect 126 38 128 66
rect 136 38 138 66
rect 146 38 148 66
rect 164 38 166 63
rect 171 38 173 63
rect 181 41 183 54
rect 194 41 196 66
rect 215 45 217 66
rect 222 45 224 66
rect 235 38 237 56
rect 36 -66 38 -41
rect 49 -54 51 -41
rect 59 -63 61 -38
rect 66 -63 68 -38
rect 84 -66 86 -38
rect 94 -66 96 -38
rect 104 -66 106 -38
rect 126 -66 128 -38
rect 136 -66 138 -38
rect 146 -66 148 -38
rect 164 -63 166 -38
rect 171 -63 173 -38
rect 181 -54 183 -41
rect 194 -66 196 -41
rect 215 -66 217 -45
rect 222 -66 224 -45
rect 235 -56 237 -38
<< polyct0 >>
rect 44 34 46 36
rect 38 24 40 26
rect 94 31 96 33
rect 104 31 106 33
rect 126 31 128 33
rect 136 31 138 33
rect 186 34 188 36
rect 233 31 235 33
rect 192 24 194 26
rect 38 -26 40 -24
rect 44 -36 46 -34
rect 94 -33 96 -31
rect 104 -33 106 -31
rect 126 -33 128 -31
rect 136 -33 138 -31
rect 192 -26 194 -24
rect 186 -36 188 -34
rect 233 -33 235 -31
<< polyct1 >>
rect 58 31 60 33
rect 77 31 79 33
rect 84 31 86 33
rect 146 31 148 33
rect 153 31 155 33
rect 172 31 174 33
rect 213 38 215 40
rect 223 31 225 33
rect 58 -33 60 -31
rect 77 -33 79 -31
rect 84 -33 86 -31
rect 146 -33 148 -31
rect 153 -33 155 -31
rect 172 -33 174 -31
rect 223 -33 225 -31
rect 213 -40 215 -38
<< ndifct0 >>
rect 41 11 43 13
rect 51 14 53 16
rect 61 22 63 24
rect 71 22 73 24
rect 71 15 73 17
rect 81 15 83 17
rect 98 8 100 10
rect 132 8 134 10
rect 159 22 161 24
rect 149 15 151 17
rect 159 15 161 17
rect 169 22 171 24
rect 220 22 222 24
rect 179 14 181 16
rect 189 11 191 13
rect 210 9 212 11
rect 229 9 231 11
rect 41 -13 43 -11
rect 51 -16 53 -14
rect 61 -24 63 -22
rect 71 -17 73 -15
rect 81 -17 83 -15
rect 71 -24 73 -22
rect 98 -10 100 -8
rect 132 -10 134 -8
rect 149 -17 151 -15
rect 159 -17 161 -15
rect 159 -24 161 -22
rect 169 -24 171 -22
rect 179 -16 181 -14
rect 189 -13 191 -11
rect 210 -11 212 -9
rect 229 -11 231 -9
rect 220 -24 222 -22
<< ndifct1 >>
rect 31 15 33 17
rect 109 15 111 17
rect 121 15 123 17
rect 199 15 201 17
rect 240 22 242 24
rect 31 -17 33 -15
rect 109 -17 111 -15
rect 121 -17 123 -15
rect 199 -17 201 -15
rect 240 -24 242 -22
<< ntiect1 >>
rect 239 65 241 67
rect 239 -67 241 -65
<< ptiect1 >>
rect 239 5 241 7
rect 239 -7 241 -5
<< pdifct0 >>
rect 42 62 44 64
rect 54 43 56 45
rect 77 62 79 64
rect 77 55 79 57
rect 89 54 91 56
rect 89 47 91 49
rect 99 62 101 64
rect 99 55 101 57
rect 131 62 133 64
rect 131 55 133 57
rect 141 54 143 56
rect 141 47 143 49
rect 153 62 155 64
rect 153 55 155 57
rect 188 62 190 64
rect 176 43 178 45
rect 210 55 212 57
rect 229 62 231 64
rect 54 -45 56 -43
rect 42 -64 44 -62
rect 77 -57 79 -55
rect 77 -64 79 -62
rect 89 -49 91 -47
rect 89 -56 91 -54
rect 99 -57 101 -55
rect 99 -64 101 -62
rect 131 -57 133 -55
rect 131 -64 133 -62
rect 141 -49 143 -47
rect 141 -56 143 -54
rect 153 -57 155 -55
rect 153 -64 155 -62
rect 176 -45 178 -43
rect 188 -64 190 -62
rect 210 -57 212 -55
rect 229 -64 231 -62
<< pdifct1 >>
rect 31 50 33 52
rect 31 43 33 45
rect 109 47 111 49
rect 109 40 111 42
rect 121 47 123 49
rect 121 40 123 42
rect 199 50 201 52
rect 199 43 201 45
rect 240 52 242 54
rect 240 45 242 47
rect 31 -45 33 -43
rect 31 -52 33 -50
rect 109 -42 111 -40
rect 109 -49 111 -47
rect 121 -42 123 -40
rect 121 -49 123 -47
rect 199 -45 201 -43
rect 199 -52 201 -50
rect 240 -47 242 -45
rect 240 -54 242 -52
<< alu0 >>
rect 40 62 42 64
rect 44 62 46 64
rect 40 61 46 62
rect 75 62 77 64
rect 79 62 81 64
rect 75 57 81 62
rect 97 62 99 64
rect 101 62 103 64
rect 75 55 77 57
rect 79 55 81 57
rect 75 54 81 55
rect 88 56 92 58
rect 88 54 89 56
rect 91 54 92 56
rect 97 57 103 62
rect 97 55 99 57
rect 101 55 103 57
rect 97 54 103 55
rect 129 62 131 64
rect 133 62 135 64
rect 129 57 135 62
rect 151 62 153 64
rect 155 62 157 64
rect 129 55 131 57
rect 133 55 135 57
rect 129 54 135 55
rect 140 56 144 58
rect 140 54 141 56
rect 143 54 144 56
rect 151 57 157 62
rect 186 62 188 64
rect 190 62 192 64
rect 186 61 192 62
rect 227 62 229 64
rect 231 62 233 64
rect 227 61 233 62
rect 151 55 153 57
rect 155 55 157 57
rect 151 54 157 55
rect 208 57 225 58
rect 208 55 210 57
rect 212 55 225 57
rect 208 54 225 55
rect 45 50 69 54
rect 88 50 92 54
rect 43 46 49 50
rect 65 49 105 50
rect 65 47 89 49
rect 91 47 105 49
rect 43 36 47 46
rect 53 45 57 47
rect 65 46 105 47
rect 53 43 54 45
rect 56 43 57 45
rect 53 42 57 43
rect 43 34 44 36
rect 46 34 47 36
rect 43 32 47 34
rect 50 38 57 42
rect 50 27 54 38
rect 93 33 97 38
rect 93 31 94 33
rect 96 31 97 33
rect 36 26 54 27
rect 36 24 38 26
rect 40 25 54 26
rect 40 24 65 25
rect 36 23 61 24
rect 50 22 61 23
rect 63 22 65 24
rect 50 21 65 22
rect 70 24 74 26
rect 70 22 71 24
rect 73 22 74 24
rect 70 17 74 22
rect 93 29 97 31
rect 101 35 105 46
rect 101 33 107 35
rect 101 31 104 33
rect 106 31 107 33
rect 101 29 107 31
rect 101 26 105 29
rect 85 22 105 26
rect 85 18 89 22
rect 49 16 71 17
rect 40 13 44 15
rect 49 14 51 16
rect 53 15 71 16
rect 73 15 74 17
rect 53 14 74 15
rect 79 17 89 18
rect 79 15 81 17
rect 83 15 89 17
rect 79 14 89 15
rect 140 50 144 54
rect 163 50 187 54
rect 127 49 167 50
rect 127 47 141 49
rect 143 47 167 49
rect 127 46 167 47
rect 127 35 131 46
rect 175 45 179 47
rect 183 46 189 50
rect 175 43 176 45
rect 178 43 179 45
rect 175 42 179 43
rect 175 38 182 42
rect 125 33 131 35
rect 125 31 126 33
rect 128 31 131 33
rect 125 29 131 31
rect 135 33 139 38
rect 135 31 136 33
rect 138 31 139 33
rect 135 29 139 31
rect 127 26 131 29
rect 127 22 147 26
rect 143 18 147 22
rect 178 27 182 38
rect 185 36 189 46
rect 185 34 186 36
rect 188 34 189 36
rect 185 32 189 34
rect 178 26 196 27
rect 158 24 162 26
rect 178 25 192 26
rect 158 22 159 24
rect 161 22 162 24
rect 143 17 153 18
rect 143 15 149 17
rect 151 15 153 17
rect 143 14 153 15
rect 158 17 162 22
rect 167 24 192 25
rect 194 24 196 26
rect 167 22 169 24
rect 171 23 196 24
rect 171 22 182 23
rect 167 21 182 22
rect 221 50 225 54
rect 221 46 236 50
rect 211 37 217 38
rect 232 33 236 46
rect 239 43 240 54
rect 232 31 233 33
rect 235 31 236 33
rect 232 25 236 31
rect 218 24 236 25
rect 218 22 220 24
rect 222 22 236 24
rect 218 21 236 22
rect 158 15 159 17
rect 161 16 183 17
rect 161 15 179 16
rect 158 14 179 15
rect 181 14 183 16
rect 49 13 74 14
rect 158 13 183 14
rect 188 13 192 15
rect 40 11 41 13
rect 43 11 44 13
rect 188 11 189 13
rect 191 11 192 13
rect 40 8 44 11
rect 96 10 102 11
rect 96 8 98 10
rect 100 8 102 10
rect 130 10 136 11
rect 130 8 132 10
rect 134 8 136 10
rect 188 8 192 11
rect 208 11 214 12
rect 208 9 210 11
rect 212 9 214 11
rect 208 8 214 9
rect 227 11 233 12
rect 227 9 229 11
rect 231 9 233 11
rect 227 8 233 9
rect 40 -11 44 -8
rect 96 -10 98 -8
rect 100 -10 102 -8
rect 96 -11 102 -10
rect 130 -10 132 -8
rect 134 -10 136 -8
rect 130 -11 136 -10
rect 188 -11 192 -8
rect 40 -13 41 -11
rect 43 -13 44 -11
rect 188 -13 189 -11
rect 191 -13 192 -11
rect 208 -9 214 -8
rect 208 -11 210 -9
rect 212 -11 214 -9
rect 208 -12 214 -11
rect 227 -9 233 -8
rect 227 -11 229 -9
rect 231 -11 233 -9
rect 227 -12 233 -11
rect 40 -15 44 -13
rect 49 -14 74 -13
rect 158 -14 183 -13
rect 49 -16 51 -14
rect 53 -15 74 -14
rect 53 -16 71 -15
rect 49 -17 71 -16
rect 73 -17 74 -15
rect 50 -22 65 -21
rect 50 -23 61 -22
rect 36 -24 61 -23
rect 63 -24 65 -22
rect 36 -26 38 -24
rect 40 -25 65 -24
rect 70 -22 74 -17
rect 79 -15 89 -14
rect 79 -17 81 -15
rect 83 -17 89 -15
rect 79 -18 89 -17
rect 70 -24 71 -22
rect 73 -24 74 -22
rect 40 -26 54 -25
rect 70 -26 74 -24
rect 36 -27 54 -26
rect 43 -34 47 -32
rect 43 -36 44 -34
rect 46 -36 47 -34
rect 43 -46 47 -36
rect 50 -38 54 -27
rect 85 -22 89 -18
rect 85 -26 105 -22
rect 101 -29 105 -26
rect 93 -31 97 -29
rect 93 -33 94 -31
rect 96 -33 97 -31
rect 93 -38 97 -33
rect 101 -31 107 -29
rect 101 -33 104 -31
rect 106 -33 107 -31
rect 101 -35 107 -33
rect 50 -42 57 -38
rect 53 -43 57 -42
rect 53 -45 54 -43
rect 56 -45 57 -43
rect 43 -50 49 -46
rect 53 -47 57 -45
rect 101 -46 105 -35
rect 65 -47 105 -46
rect 65 -49 89 -47
rect 91 -49 105 -47
rect 65 -50 105 -49
rect 45 -54 69 -50
rect 88 -54 92 -50
rect 143 -15 153 -14
rect 143 -17 149 -15
rect 151 -17 153 -15
rect 143 -18 153 -17
rect 158 -15 179 -14
rect 158 -17 159 -15
rect 161 -16 179 -15
rect 181 -16 183 -14
rect 188 -15 192 -13
rect 161 -17 183 -16
rect 143 -22 147 -18
rect 127 -26 147 -22
rect 127 -29 131 -26
rect 125 -31 131 -29
rect 125 -33 126 -31
rect 128 -33 131 -31
rect 125 -35 131 -33
rect 127 -46 131 -35
rect 135 -31 139 -29
rect 158 -22 162 -17
rect 158 -24 159 -22
rect 161 -24 162 -22
rect 158 -26 162 -24
rect 167 -22 182 -21
rect 167 -24 169 -22
rect 171 -23 182 -22
rect 171 -24 196 -23
rect 167 -25 192 -24
rect 178 -26 192 -25
rect 194 -26 196 -24
rect 178 -27 196 -26
rect 135 -33 136 -31
rect 138 -33 139 -31
rect 135 -38 139 -33
rect 178 -38 182 -27
rect 175 -42 182 -38
rect 185 -34 189 -32
rect 185 -36 186 -34
rect 188 -36 189 -34
rect 175 -43 179 -42
rect 175 -45 176 -43
rect 178 -45 179 -43
rect 127 -47 167 -46
rect 175 -47 179 -45
rect 185 -46 189 -36
rect 218 -22 236 -21
rect 218 -24 220 -22
rect 222 -24 236 -22
rect 218 -25 236 -24
rect 232 -31 236 -25
rect 232 -33 233 -31
rect 235 -33 236 -31
rect 211 -38 217 -37
rect 127 -49 141 -47
rect 143 -49 167 -47
rect 127 -50 167 -49
rect 183 -50 189 -46
rect 140 -54 144 -50
rect 163 -54 187 -50
rect 232 -46 236 -33
rect 221 -50 236 -46
rect 221 -54 225 -50
rect 239 -54 240 -43
rect 75 -55 81 -54
rect 75 -57 77 -55
rect 79 -57 81 -55
rect 40 -62 46 -61
rect 40 -64 42 -62
rect 44 -64 46 -62
rect 75 -62 81 -57
rect 88 -56 89 -54
rect 91 -56 92 -54
rect 88 -58 92 -56
rect 97 -55 103 -54
rect 97 -57 99 -55
rect 101 -57 103 -55
rect 75 -64 77 -62
rect 79 -64 81 -62
rect 97 -62 103 -57
rect 97 -64 99 -62
rect 101 -64 103 -62
rect 129 -55 135 -54
rect 129 -57 131 -55
rect 133 -57 135 -55
rect 129 -62 135 -57
rect 140 -56 141 -54
rect 143 -56 144 -54
rect 140 -58 144 -56
rect 151 -55 157 -54
rect 151 -57 153 -55
rect 155 -57 157 -55
rect 129 -64 131 -62
rect 133 -64 135 -62
rect 151 -62 157 -57
rect 208 -55 225 -54
rect 208 -57 210 -55
rect 212 -57 225 -55
rect 208 -58 225 -57
rect 151 -64 153 -62
rect 155 -64 157 -62
rect 186 -62 192 -61
rect 186 -64 188 -62
rect 190 -64 192 -62
rect 227 -62 233 -61
rect 227 -64 229 -62
rect 231 -64 233 -62
<< via1 >>
rect 30 23 32 25
rect 111 31 113 33
rect 121 44 123 46
rect 152 23 154 25
rect 209 44 211 46
rect 209 31 211 33
rect 241 27 243 29
rect 30 -25 32 -23
rect 111 -33 113 -31
rect 152 -25 154 -23
rect 121 -46 123 -44
rect 169 -38 171 -36
rect 209 -27 211 -25
rect 209 -46 211 -44
<< via2 >>
rect 245 27 247 29
rect 245 -38 247 -36
<< labels >>
rlabel alu1 75 4 75 4 1 gnd
rlabel alu1 157 4 157 4 1 gnd
rlabel alu1 154 40 154 40 1 cin
rlabel alu1 242 -38 242 -38 5 cout
rlabel alu1 157 -4 157 -4 5 gnd
rlabel alu1 75 -4 75 -4 5 gnd
rlabel alu1 79 40 79 40 1 b_0
rlabel alu1 87 32 87 32 1 a_0
rlabel alu1 87 -32 87 -32 1 a_1
rlabel alu1 79 -40 79 -40 1 b_1
rlabel alu1 201 -32 201 -32 1 s_1
rlabel alu1 201 37 201 37 1 s_0
rlabel alu1 180 68 180 68 1 Vdd
rlabel alu1 206 68 206 68 1 Vdd
rlabel alu1 116 68 116 68 1 Vdd
rlabel alu1 51 68 51 68 1 vdd
rlabel alu1 51 -69 51 -69 1 Vdd
rlabel alu1 116 -68 116 -68 1 Vdd
rlabel alu1 207 -68 207 -68 1 Vdd
rlabel alu1 181 -68 181 -68 1 Vdd
<< end >>
