magic
tech scmos
timestamp 1520963264
<< nwell >>
rect -16 -3 17 18
<< polysilicon >>
rect -13 9 -11 11
rect -2 9 0 11
rect 7 9 9 11
rect -13 -9 -11 -3
rect -2 -9 0 -3
rect 7 -9 9 -3
rect -12 -13 -11 -9
rect -1 -13 0 -9
rect -13 -21 -11 -13
rect -2 -21 0 -13
rect 7 -24 9 -13
rect -13 -29 -11 -27
rect -2 -29 0 -27
rect 7 -29 9 -27
<< ndiffusion >>
rect -16 -22 -13 -21
rect -14 -26 -13 -22
rect -16 -27 -13 -26
rect -11 -27 -2 -21
rect 0 -22 6 -21
rect 0 -26 1 -22
rect 5 -24 6 -22
rect 5 -26 7 -24
rect 0 -27 7 -26
rect 9 -27 12 -24
rect 16 -27 17 -24
<< pdiffusion >>
rect -16 5 -13 9
rect -15 1 -13 5
rect -16 -3 -13 1
rect -11 5 -2 9
rect -11 1 -8 5
rect -4 1 -2 5
rect -11 -3 -2 1
rect 0 5 7 9
rect 0 1 2 5
rect 6 1 7 5
rect 0 -3 7 1
rect 9 5 17 9
rect 9 1 11 5
rect 15 1 17 5
rect 9 -3 17 1
<< metal1 >>
rect -18 17 17 18
rect -18 15 12 17
rect -8 5 -5 15
rect 16 15 17 17
rect -18 -3 -15 1
rect 2 -3 5 1
rect -18 -6 5 -3
rect 12 -16 15 1
rect -18 -19 15 -16
rect -18 -22 -15 -19
rect 2 -31 5 -26
rect 12 -23 15 -19
rect -18 -34 17 -31
<< ntransistor >>
rect -13 -27 -11 -21
rect -2 -27 0 -21
rect 7 -27 9 -24
<< ptransistor >>
rect -13 -3 -11 9
rect -2 -3 0 9
rect 7 -3 9 9
<< polycontact >>
rect -16 -13 -12 -9
rect -5 -13 -1 -9
rect 5 -13 9 -9
<< ndcontact >>
rect -18 -26 -14 -22
rect 1 -26 5 -22
rect 12 -27 16 -23
<< pdcontact >>
rect -19 1 -15 5
rect -8 1 -4 5
rect 2 1 6 5
rect 11 1 15 5
<< nsubstratencontact >>
rect 12 13 16 17
<< labels >>
rlabel metal1 -11 17 -11 17 5 vdd
rlabel polycontact -15 -11 -15 -11 3 B
rlabel polycontact -3 -11 -3 -11 1 C
rlabel polycontact 7 -11 7 -11 1 A
rlabel ndiffusion -7 -24 -7 -24 1 n1
rlabel metal1 -2 -33 -2 -33 1 gnd
rlabel metal1 14 -11 14 -11 1 out
rlabel pdcontact 4 3 4 3 1 n2
<< end >>
