* SPICE3 file created from (UNNAMED).ext - technology: scmos

.include /home/vlsilab/UG_students_2018/t14y_tsmc_025_level3.txt


M1000 out in vdd vdd cmosp w=3u l=2u
+  ad=19p pd=18u as=19p ps=18u
M1001 out in gnd Gnd cmosn w=3u l=2u
+  ad=19p pd=18u as=19p ps=18u

C0 in vdd 2.15fF
C1 gnd Gnd 3.81fF
C2 in Gnd 4.52fF
C3 vdd Gnd 2.82fF

v_dd vdd 0 5
gd gnd 0 0
gd Gnd 0 0 

v_in in 0 PULSE(0 5 0 0.1n 0.1n 5n 10n)



.control
tran 0.01n 40n
run
plot (in) (out)


plot vdd*(-v_dd#branch)


meas tran yavg AVG i(v_dd) from=0ns to=10ns

.endc

print yavg
.end


