* SPICE3 file created from nand2.ext - technology: scmos

.option scale=1u

M1000 Out InB Vdd Vdd pfet w=3 l=2
+  ad=22 pd=20 as=50 ps=44
M1001 Vdd InA Out Vdd pfet w=3 l=2
+  ad=0 pd=0 as=0 ps=0
M1002 a_4_0# InB Gnd Gnd nfet w=3 l=2
+  ad=18 pd=18 as=25 ps=22
M1003 Out InA a_4_0# Gnd nfet w=3 l=2
+  ad=25 pd=22 as=0 ps=0
C0 Gnd Gnd 3.95fF
C1 InA Gnd 6.14fF
C2 InB Gnd 3.81fF
