magic
tech scmos
timestamp 1520355758
<< nwell >>
rect -4 24 8 25
rect -7 4 8 24
<< polysilicon >>
rect -2 13 2 16
rect -2 2 2 9
rect -1 -4 1 -2
rect -1 -10 1 -8
<< ndiffusion >>
rect -5 -8 -1 -4
rect 1 -8 5 -4
<< pdiffusion >>
rect -5 9 -2 13
rect 2 9 5 13
<< metal1 >>
rect -8 30 8 33
rect -8 26 -5 30
rect -9 22 -8 26
rect -9 14 -6 22
rect 6 -4 9 9
rect -8 -12 -5 -8
rect -8 -15 9 -12
<< ntransistor >>
rect -1 -8 1 -4
<< ptransistor >>
rect -2 9 2 13
<< polycontact >>
rect -2 -2 2 2
<< ndcontact >>
rect -9 -8 -5 -4
rect 5 -8 9 -4
<< pdcontact >>
rect -9 9 -5 14
rect 5 9 9 14
<< nsubstratencontact >>
rect -8 22 -4 26
<< labels >>
rlabel polycontact 0 0 0 0 1 in
rlabel metal1 0 -14 0 -14 1 gnd
rlabel metal1 8 0 8 0 7 out
rlabel metal1 0 31 0 31 5 vdd
<< end >>
