magic
tech scmos
timestamp 1553838827
<< rotate >>
rect 75 12 86 14
rect 52 8 54 10
rect 75 5 89 12
rect 78 3 89 5
rect 75 -132 86 -130
rect 52 -136 54 -134
rect 75 -139 89 -132
rect 78 -141 89 -139
<< ab >>
rect 5 135 182 149
rect 5 131 7 135
rect 9 131 179 135
rect 181 131 182 135
rect 5 23 182 131
rect 5 19 7 23
rect 9 19 179 23
rect 181 19 182 23
rect 5 -9 182 19
rect 5 -13 7 -9
rect 9 -13 179 -9
rect 181 -13 182 -9
rect 5 -121 182 -13
rect 5 -125 7 -121
rect 9 -125 179 -121
rect 181 -125 182 -121
rect 5 -139 182 -125
rect 184 38 225 149
rect 184 35 226 38
rect 184 -106 225 35
rect 184 -109 226 -106
rect 184 -139 225 -109
<< nwell >>
rect 0 109 228 154
rect 0 -35 228 45
rect 0 -144 228 -99
<< pwell >>
rect 0 45 228 109
rect 0 -99 228 -35
<< poly >>
rect 14 143 16 147
rect 37 140 39 145
rect 44 140 46 145
rect 62 143 64 147
rect 72 143 74 147
rect 82 143 84 147
rect 104 143 106 147
rect 114 143 116 147
rect 124 143 126 147
rect 27 131 29 136
rect 14 105 16 118
rect 27 115 29 118
rect 142 140 144 145
rect 149 140 151 145
rect 172 143 174 147
rect 193 143 195 147
rect 200 143 202 147
rect 159 131 161 136
rect 213 133 215 138
rect 193 119 195 122
rect 159 115 161 118
rect 20 113 29 115
rect 20 111 22 113
rect 24 111 26 113
rect 37 112 39 115
rect 44 112 46 115
rect 62 112 64 115
rect 72 112 74 115
rect 82 112 84 115
rect 104 112 106 115
rect 114 112 116 115
rect 124 112 126 115
rect 142 112 144 115
rect 149 112 151 115
rect 159 113 168 115
rect 20 109 26 111
rect 14 103 20 105
rect 14 101 16 103
rect 18 101 20 103
rect 14 99 20 101
rect 14 96 16 99
rect 24 96 26 109
rect 34 110 40 112
rect 34 108 36 110
rect 38 108 40 110
rect 34 106 40 108
rect 44 110 66 112
rect 44 108 55 110
rect 57 108 62 110
rect 64 108 66 110
rect 44 106 66 108
rect 70 110 76 112
rect 70 108 72 110
rect 74 108 76 110
rect 70 106 76 108
rect 80 110 86 112
rect 80 108 82 110
rect 84 108 86 110
rect 80 106 86 108
rect 102 110 108 112
rect 102 108 104 110
rect 106 108 108 110
rect 102 106 108 108
rect 112 110 118 112
rect 112 108 114 110
rect 116 108 118 110
rect 112 106 118 108
rect 122 110 144 112
rect 122 108 124 110
rect 126 108 131 110
rect 133 108 144 110
rect 122 106 144 108
rect 148 110 154 112
rect 148 108 150 110
rect 152 108 154 110
rect 148 106 154 108
rect 34 103 36 106
rect 44 103 46 106
rect 64 103 66 106
rect 71 103 73 106
rect 14 79 16 83
rect 24 81 26 86
rect 34 84 36 89
rect 44 84 46 89
rect 82 97 84 106
rect 104 97 106 106
rect 115 103 117 106
rect 122 103 124 106
rect 142 103 144 106
rect 152 103 154 106
rect 162 111 164 113
rect 166 111 168 113
rect 162 109 168 111
rect 162 96 164 109
rect 172 105 174 118
rect 189 117 195 119
rect 189 115 191 117
rect 193 115 195 117
rect 189 113 195 115
rect 168 103 174 105
rect 193 103 195 113
rect 200 112 202 122
rect 213 112 215 115
rect 199 110 205 112
rect 199 108 201 110
rect 203 108 205 110
rect 199 106 205 108
rect 209 110 215 112
rect 209 108 211 110
rect 213 108 215 110
rect 209 106 215 108
rect 203 103 205 106
rect 213 103 215 106
rect 168 101 170 103
rect 172 101 174 103
rect 168 99 174 101
rect 172 96 174 99
rect 142 84 144 89
rect 152 84 154 89
rect 64 79 66 83
rect 71 79 73 83
rect 82 79 84 83
rect 104 79 106 83
rect 115 79 117 83
rect 122 79 124 83
rect 162 81 164 86
rect 193 92 195 97
rect 203 92 205 97
rect 213 89 215 94
rect 172 79 174 83
rect 14 71 16 75
rect 24 68 26 73
rect 64 71 66 75
rect 71 71 73 75
rect 82 71 84 75
rect 104 71 106 75
rect 115 71 117 75
rect 122 71 124 75
rect 34 65 36 70
rect 44 65 46 70
rect 14 55 16 58
rect 14 53 20 55
rect 14 51 16 53
rect 18 51 20 53
rect 14 49 20 51
rect 14 36 16 49
rect 24 45 26 58
rect 20 43 26 45
rect 20 41 22 43
rect 24 41 26 43
rect 34 48 36 51
rect 44 48 46 51
rect 64 48 66 51
rect 71 48 73 51
rect 82 48 84 57
rect 104 48 106 57
rect 142 65 144 70
rect 152 65 154 70
rect 162 68 164 73
rect 172 71 174 75
rect 115 48 117 51
rect 122 48 124 51
rect 142 48 144 51
rect 152 48 154 51
rect 34 46 40 48
rect 34 44 36 46
rect 38 44 40 46
rect 34 42 40 44
rect 44 46 66 48
rect 44 44 55 46
rect 57 44 62 46
rect 64 44 66 46
rect 44 42 66 44
rect 70 46 76 48
rect 70 44 72 46
rect 74 44 76 46
rect 70 42 76 44
rect 80 46 86 48
rect 80 44 82 46
rect 84 44 86 46
rect 80 42 86 44
rect 102 46 108 48
rect 102 44 104 46
rect 106 44 108 46
rect 102 42 108 44
rect 112 46 118 48
rect 112 44 114 46
rect 116 44 118 46
rect 112 42 118 44
rect 122 46 144 48
rect 122 44 124 46
rect 126 44 131 46
rect 133 44 144 46
rect 122 42 144 44
rect 148 46 154 48
rect 148 44 150 46
rect 152 44 154 46
rect 148 42 154 44
rect 162 45 164 58
rect 172 55 174 58
rect 168 53 174 55
rect 168 51 170 53
rect 172 51 174 53
rect 193 57 195 62
rect 203 57 205 62
rect 213 60 215 65
rect 168 49 174 51
rect 162 43 168 45
rect 20 39 29 41
rect 37 39 39 42
rect 44 39 46 42
rect 62 39 64 42
rect 72 39 74 42
rect 82 39 84 42
rect 104 39 106 42
rect 114 39 116 42
rect 124 39 126 42
rect 142 39 144 42
rect 149 39 151 42
rect 162 41 164 43
rect 166 41 168 43
rect 159 39 168 41
rect 27 36 29 39
rect 27 18 29 23
rect 14 7 16 11
rect 37 9 39 14
rect 44 9 46 14
rect 159 36 161 39
rect 172 36 174 49
rect 193 41 195 51
rect 203 48 205 51
rect 213 48 215 51
rect 199 46 205 48
rect 199 44 201 46
rect 203 44 205 46
rect 199 42 205 44
rect 209 46 215 48
rect 209 44 211 46
rect 213 44 215 46
rect 209 42 215 44
rect 189 39 195 41
rect 189 37 191 39
rect 193 37 195 39
rect 159 18 161 23
rect 62 7 64 11
rect 72 7 74 11
rect 82 7 84 11
rect 104 7 106 11
rect 114 7 116 11
rect 124 7 126 11
rect 142 9 144 14
rect 149 9 151 14
rect 189 35 195 37
rect 193 32 195 35
rect 200 32 202 42
rect 213 39 215 42
rect 213 16 215 21
rect 172 7 174 11
rect 193 7 195 11
rect 200 7 202 11
rect 14 -1 16 3
rect 37 -4 39 1
rect 44 -4 46 1
rect 62 -1 64 3
rect 72 -1 74 3
rect 82 -1 84 3
rect 104 -1 106 3
rect 114 -1 116 3
rect 124 -1 126 3
rect 27 -13 29 -8
rect 14 -39 16 -26
rect 27 -29 29 -26
rect 142 -4 144 1
rect 149 -4 151 1
rect 172 -1 174 3
rect 193 -1 195 3
rect 200 -1 202 3
rect 159 -13 161 -8
rect 213 -11 215 -6
rect 193 -25 195 -22
rect 159 -29 161 -26
rect 20 -31 29 -29
rect 20 -33 22 -31
rect 24 -33 26 -31
rect 37 -32 39 -29
rect 44 -32 46 -29
rect 62 -32 64 -29
rect 72 -32 74 -29
rect 82 -32 84 -29
rect 104 -32 106 -29
rect 114 -32 116 -29
rect 124 -32 126 -29
rect 142 -32 144 -29
rect 149 -32 151 -29
rect 159 -31 168 -29
rect 20 -35 26 -33
rect 14 -41 20 -39
rect 14 -43 16 -41
rect 18 -43 20 -41
rect 14 -45 20 -43
rect 14 -48 16 -45
rect 24 -48 26 -35
rect 34 -34 40 -32
rect 34 -36 36 -34
rect 38 -36 40 -34
rect 34 -38 40 -36
rect 44 -34 66 -32
rect 44 -36 55 -34
rect 57 -36 62 -34
rect 64 -36 66 -34
rect 44 -38 66 -36
rect 70 -34 76 -32
rect 70 -36 72 -34
rect 74 -36 76 -34
rect 70 -38 76 -36
rect 80 -34 86 -32
rect 80 -36 82 -34
rect 84 -36 86 -34
rect 80 -38 86 -36
rect 102 -34 108 -32
rect 102 -36 104 -34
rect 106 -36 108 -34
rect 102 -38 108 -36
rect 112 -34 118 -32
rect 112 -36 114 -34
rect 116 -36 118 -34
rect 112 -38 118 -36
rect 122 -34 144 -32
rect 122 -36 124 -34
rect 126 -36 131 -34
rect 133 -36 144 -34
rect 122 -38 144 -36
rect 148 -34 154 -32
rect 148 -36 150 -34
rect 152 -36 154 -34
rect 148 -38 154 -36
rect 34 -41 36 -38
rect 44 -41 46 -38
rect 64 -41 66 -38
rect 71 -41 73 -38
rect 14 -65 16 -61
rect 24 -63 26 -58
rect 34 -60 36 -55
rect 44 -60 46 -55
rect 82 -47 84 -38
rect 104 -47 106 -38
rect 115 -41 117 -38
rect 122 -41 124 -38
rect 142 -41 144 -38
rect 152 -41 154 -38
rect 162 -33 164 -31
rect 166 -33 168 -31
rect 162 -35 168 -33
rect 162 -48 164 -35
rect 172 -39 174 -26
rect 189 -27 195 -25
rect 189 -29 191 -27
rect 193 -29 195 -27
rect 189 -31 195 -29
rect 168 -41 174 -39
rect 193 -41 195 -31
rect 200 -32 202 -22
rect 213 -32 215 -29
rect 199 -34 205 -32
rect 199 -36 201 -34
rect 203 -36 205 -34
rect 199 -38 205 -36
rect 209 -34 215 -32
rect 209 -36 211 -34
rect 213 -36 215 -34
rect 209 -38 215 -36
rect 203 -41 205 -38
rect 213 -41 215 -38
rect 168 -43 170 -41
rect 172 -43 174 -41
rect 168 -45 174 -43
rect 172 -48 174 -45
rect 142 -60 144 -55
rect 152 -60 154 -55
rect 64 -65 66 -61
rect 71 -65 73 -61
rect 82 -65 84 -61
rect 104 -65 106 -61
rect 115 -65 117 -61
rect 122 -65 124 -61
rect 162 -63 164 -58
rect 193 -52 195 -47
rect 203 -52 205 -47
rect 213 -55 215 -50
rect 172 -65 174 -61
rect 14 -73 16 -69
rect 24 -76 26 -71
rect 64 -73 66 -69
rect 71 -73 73 -69
rect 82 -73 84 -69
rect 104 -73 106 -69
rect 115 -73 117 -69
rect 122 -73 124 -69
rect 34 -79 36 -74
rect 44 -79 46 -74
rect 14 -89 16 -86
rect 14 -91 20 -89
rect 14 -93 16 -91
rect 18 -93 20 -91
rect 14 -95 20 -93
rect 14 -108 16 -95
rect 24 -99 26 -86
rect 20 -101 26 -99
rect 20 -103 22 -101
rect 24 -103 26 -101
rect 34 -96 36 -93
rect 44 -96 46 -93
rect 64 -96 66 -93
rect 71 -96 73 -93
rect 82 -96 84 -87
rect 104 -96 106 -87
rect 142 -79 144 -74
rect 152 -79 154 -74
rect 162 -76 164 -71
rect 172 -73 174 -69
rect 115 -96 117 -93
rect 122 -96 124 -93
rect 142 -96 144 -93
rect 152 -96 154 -93
rect 34 -98 40 -96
rect 34 -100 36 -98
rect 38 -100 40 -98
rect 34 -102 40 -100
rect 44 -98 66 -96
rect 44 -100 55 -98
rect 57 -100 62 -98
rect 64 -100 66 -98
rect 44 -102 66 -100
rect 70 -98 76 -96
rect 70 -100 72 -98
rect 74 -100 76 -98
rect 70 -102 76 -100
rect 80 -98 86 -96
rect 80 -100 82 -98
rect 84 -100 86 -98
rect 80 -102 86 -100
rect 102 -98 108 -96
rect 102 -100 104 -98
rect 106 -100 108 -98
rect 102 -102 108 -100
rect 112 -98 118 -96
rect 112 -100 114 -98
rect 116 -100 118 -98
rect 112 -102 118 -100
rect 122 -98 144 -96
rect 122 -100 124 -98
rect 126 -100 131 -98
rect 133 -100 144 -98
rect 122 -102 144 -100
rect 148 -98 154 -96
rect 148 -100 150 -98
rect 152 -100 154 -98
rect 148 -102 154 -100
rect 162 -99 164 -86
rect 172 -89 174 -86
rect 168 -91 174 -89
rect 168 -93 170 -91
rect 172 -93 174 -91
rect 193 -87 195 -82
rect 203 -87 205 -82
rect 213 -84 215 -79
rect 168 -95 174 -93
rect 162 -101 168 -99
rect 20 -105 29 -103
rect 37 -105 39 -102
rect 44 -105 46 -102
rect 62 -105 64 -102
rect 72 -105 74 -102
rect 82 -105 84 -102
rect 104 -105 106 -102
rect 114 -105 116 -102
rect 124 -105 126 -102
rect 142 -105 144 -102
rect 149 -105 151 -102
rect 162 -103 164 -101
rect 166 -103 168 -101
rect 159 -105 168 -103
rect 27 -108 29 -105
rect 27 -126 29 -121
rect 14 -137 16 -133
rect 37 -135 39 -130
rect 44 -135 46 -130
rect 159 -108 161 -105
rect 172 -108 174 -95
rect 193 -103 195 -93
rect 203 -96 205 -93
rect 213 -96 215 -93
rect 199 -98 205 -96
rect 199 -100 201 -98
rect 203 -100 205 -98
rect 199 -102 205 -100
rect 209 -98 215 -96
rect 209 -100 211 -98
rect 213 -100 215 -98
rect 209 -102 215 -100
rect 189 -105 195 -103
rect 189 -107 191 -105
rect 193 -107 195 -105
rect 159 -126 161 -121
rect 62 -137 64 -133
rect 72 -137 74 -133
rect 82 -137 84 -133
rect 104 -137 106 -133
rect 114 -137 116 -133
rect 124 -137 126 -133
rect 142 -135 144 -130
rect 149 -135 151 -130
rect 189 -109 195 -107
rect 193 -112 195 -109
rect 200 -112 202 -102
rect 213 -105 215 -102
rect 213 -128 215 -123
rect 172 -137 174 -133
rect 193 -137 195 -133
rect 200 -137 202 -133
<< ndif >>
rect 29 96 34 103
rect 7 94 14 96
rect 7 92 9 94
rect 11 92 14 94
rect 7 90 14 92
rect 9 83 14 90
rect 16 90 24 96
rect 16 88 19 90
rect 21 88 24 90
rect 16 86 24 88
rect 26 93 34 96
rect 26 91 29 93
rect 31 91 34 93
rect 26 89 34 91
rect 36 101 44 103
rect 36 99 39 101
rect 41 99 44 101
rect 36 89 44 99
rect 46 101 53 103
rect 46 99 49 101
rect 51 99 53 101
rect 46 94 53 99
rect 59 96 64 103
rect 46 92 49 94
rect 51 92 53 94
rect 46 89 53 92
rect 57 94 64 96
rect 57 92 59 94
rect 61 92 64 94
rect 57 90 64 92
rect 26 86 31 89
rect 16 83 21 86
rect 59 83 64 90
rect 66 83 71 103
rect 73 97 80 103
rect 108 97 115 103
rect 73 87 82 97
rect 73 85 76 87
rect 78 85 82 87
rect 73 83 82 85
rect 84 94 91 97
rect 84 92 87 94
rect 89 92 91 94
rect 84 90 91 92
rect 97 94 104 97
rect 97 92 99 94
rect 101 92 104 94
rect 97 90 104 92
rect 84 83 89 90
rect 99 83 104 90
rect 106 87 115 97
rect 106 85 110 87
rect 112 85 115 87
rect 106 83 115 85
rect 117 83 122 103
rect 124 96 129 103
rect 135 101 142 103
rect 135 99 137 101
rect 139 99 142 101
rect 124 94 131 96
rect 124 92 127 94
rect 129 92 131 94
rect 124 90 131 92
rect 135 94 142 99
rect 135 92 137 94
rect 139 92 142 94
rect 124 83 129 90
rect 135 89 142 92
rect 144 101 152 103
rect 144 99 147 101
rect 149 99 152 101
rect 144 89 152 99
rect 154 96 159 103
rect 186 97 193 103
rect 195 101 203 103
rect 195 99 198 101
rect 200 99 203 101
rect 195 97 203 99
rect 205 97 213 103
rect 154 93 162 96
rect 154 91 157 93
rect 159 91 162 93
rect 154 89 162 91
rect 157 86 162 89
rect 164 90 172 96
rect 164 88 167 90
rect 169 88 172 90
rect 164 86 172 88
rect 167 83 172 86
rect 174 94 181 96
rect 174 92 177 94
rect 179 92 181 94
rect 174 90 181 92
rect 186 90 191 97
rect 207 94 213 97
rect 215 101 222 103
rect 215 99 218 101
rect 220 99 222 101
rect 215 97 222 99
rect 215 94 220 97
rect 207 90 211 94
rect 174 83 179 90
rect 186 88 192 90
rect 186 86 188 88
rect 190 86 192 88
rect 186 84 192 86
rect 205 88 211 90
rect 205 86 207 88
rect 209 86 211 88
rect 205 84 211 86
rect 9 64 14 71
rect 7 62 14 64
rect 7 60 9 62
rect 11 60 14 62
rect 7 58 14 60
rect 16 68 21 71
rect 16 66 24 68
rect 16 64 19 66
rect 21 64 24 66
rect 16 58 24 64
rect 26 65 31 68
rect 26 63 34 65
rect 26 61 29 63
rect 31 61 34 63
rect 26 58 34 61
rect 29 51 34 58
rect 36 55 44 65
rect 36 53 39 55
rect 41 53 44 55
rect 36 51 44 53
rect 46 62 53 65
rect 59 64 64 71
rect 46 60 49 62
rect 51 60 53 62
rect 46 55 53 60
rect 57 62 64 64
rect 57 60 59 62
rect 61 60 64 62
rect 57 58 64 60
rect 46 53 49 55
rect 51 53 53 55
rect 46 51 53 53
rect 59 51 64 58
rect 66 51 71 71
rect 73 69 82 71
rect 73 67 76 69
rect 78 67 82 69
rect 73 57 82 67
rect 84 64 89 71
rect 99 64 104 71
rect 84 62 91 64
rect 84 60 87 62
rect 89 60 91 62
rect 84 57 91 60
rect 97 62 104 64
rect 97 60 99 62
rect 101 60 104 62
rect 97 57 104 60
rect 106 69 115 71
rect 106 67 110 69
rect 112 67 115 69
rect 106 57 115 67
rect 73 51 80 57
rect 108 51 115 57
rect 117 51 122 71
rect 124 64 129 71
rect 167 68 172 71
rect 157 65 162 68
rect 124 62 131 64
rect 124 60 127 62
rect 129 60 131 62
rect 124 58 131 60
rect 135 62 142 65
rect 135 60 137 62
rect 139 60 142 62
rect 124 51 129 58
rect 135 55 142 60
rect 135 53 137 55
rect 139 53 142 55
rect 135 51 142 53
rect 144 55 152 65
rect 144 53 147 55
rect 149 53 152 55
rect 144 51 152 53
rect 154 63 162 65
rect 154 61 157 63
rect 159 61 162 63
rect 154 58 162 61
rect 164 66 172 68
rect 164 64 167 66
rect 169 64 172 66
rect 164 58 172 64
rect 174 64 179 71
rect 186 68 192 70
rect 186 66 188 68
rect 190 66 192 68
rect 186 64 192 66
rect 205 68 211 70
rect 205 66 207 68
rect 209 66 211 68
rect 205 64 211 66
rect 174 62 181 64
rect 174 60 177 62
rect 179 60 181 62
rect 174 58 181 60
rect 154 51 159 58
rect 186 57 191 64
rect 207 60 211 64
rect 207 57 213 60
rect 186 51 193 57
rect 195 55 203 57
rect 195 53 198 55
rect 200 53 203 55
rect 195 51 203 53
rect 205 51 213 57
rect 215 57 220 60
rect 215 55 222 57
rect 215 53 218 55
rect 220 53 222 55
rect 215 51 222 53
rect 29 -48 34 -41
rect 7 -50 14 -48
rect 7 -52 9 -50
rect 11 -52 14 -50
rect 7 -54 14 -52
rect 9 -61 14 -54
rect 16 -54 24 -48
rect 16 -56 19 -54
rect 21 -56 24 -54
rect 16 -58 24 -56
rect 26 -51 34 -48
rect 26 -53 29 -51
rect 31 -53 34 -51
rect 26 -55 34 -53
rect 36 -43 44 -41
rect 36 -45 39 -43
rect 41 -45 44 -43
rect 36 -55 44 -45
rect 46 -43 53 -41
rect 46 -45 49 -43
rect 51 -45 53 -43
rect 46 -50 53 -45
rect 59 -48 64 -41
rect 46 -52 49 -50
rect 51 -52 53 -50
rect 46 -55 53 -52
rect 57 -50 64 -48
rect 57 -52 59 -50
rect 61 -52 64 -50
rect 57 -54 64 -52
rect 26 -58 31 -55
rect 16 -61 21 -58
rect 59 -61 64 -54
rect 66 -61 71 -41
rect 73 -47 80 -41
rect 108 -47 115 -41
rect 73 -57 82 -47
rect 73 -59 76 -57
rect 78 -59 82 -57
rect 73 -61 82 -59
rect 84 -50 91 -47
rect 84 -52 87 -50
rect 89 -52 91 -50
rect 84 -54 91 -52
rect 97 -50 104 -47
rect 97 -52 99 -50
rect 101 -52 104 -50
rect 97 -54 104 -52
rect 84 -61 89 -54
rect 99 -61 104 -54
rect 106 -57 115 -47
rect 106 -59 110 -57
rect 112 -59 115 -57
rect 106 -61 115 -59
rect 117 -61 122 -41
rect 124 -48 129 -41
rect 135 -43 142 -41
rect 135 -45 137 -43
rect 139 -45 142 -43
rect 124 -50 131 -48
rect 124 -52 127 -50
rect 129 -52 131 -50
rect 124 -54 131 -52
rect 135 -50 142 -45
rect 135 -52 137 -50
rect 139 -52 142 -50
rect 124 -61 129 -54
rect 135 -55 142 -52
rect 144 -43 152 -41
rect 144 -45 147 -43
rect 149 -45 152 -43
rect 144 -55 152 -45
rect 154 -48 159 -41
rect 186 -47 193 -41
rect 195 -43 203 -41
rect 195 -45 198 -43
rect 200 -45 203 -43
rect 195 -47 203 -45
rect 205 -47 213 -41
rect 154 -51 162 -48
rect 154 -53 157 -51
rect 159 -53 162 -51
rect 154 -55 162 -53
rect 157 -58 162 -55
rect 164 -54 172 -48
rect 164 -56 167 -54
rect 169 -56 172 -54
rect 164 -58 172 -56
rect 167 -61 172 -58
rect 174 -50 181 -48
rect 174 -52 177 -50
rect 179 -52 181 -50
rect 174 -54 181 -52
rect 186 -54 191 -47
rect 207 -50 213 -47
rect 215 -43 222 -41
rect 215 -45 218 -43
rect 220 -45 222 -43
rect 215 -47 222 -45
rect 215 -50 220 -47
rect 207 -54 211 -50
rect 174 -61 179 -54
rect 186 -56 192 -54
rect 186 -58 188 -56
rect 190 -58 192 -56
rect 186 -60 192 -58
rect 205 -56 211 -54
rect 205 -58 207 -56
rect 209 -58 211 -56
rect 205 -60 211 -58
rect 9 -80 14 -73
rect 7 -82 14 -80
rect 7 -84 9 -82
rect 11 -84 14 -82
rect 7 -86 14 -84
rect 16 -76 21 -73
rect 16 -78 24 -76
rect 16 -80 19 -78
rect 21 -80 24 -78
rect 16 -86 24 -80
rect 26 -79 31 -76
rect 26 -81 34 -79
rect 26 -83 29 -81
rect 31 -83 34 -81
rect 26 -86 34 -83
rect 29 -93 34 -86
rect 36 -89 44 -79
rect 36 -91 39 -89
rect 41 -91 44 -89
rect 36 -93 44 -91
rect 46 -82 53 -79
rect 59 -80 64 -73
rect 46 -84 49 -82
rect 51 -84 53 -82
rect 46 -89 53 -84
rect 57 -82 64 -80
rect 57 -84 59 -82
rect 61 -84 64 -82
rect 57 -86 64 -84
rect 46 -91 49 -89
rect 51 -91 53 -89
rect 46 -93 53 -91
rect 59 -93 64 -86
rect 66 -93 71 -73
rect 73 -75 82 -73
rect 73 -77 76 -75
rect 78 -77 82 -75
rect 73 -87 82 -77
rect 84 -80 89 -73
rect 99 -80 104 -73
rect 84 -82 91 -80
rect 84 -84 87 -82
rect 89 -84 91 -82
rect 84 -87 91 -84
rect 97 -82 104 -80
rect 97 -84 99 -82
rect 101 -84 104 -82
rect 97 -87 104 -84
rect 106 -75 115 -73
rect 106 -77 110 -75
rect 112 -77 115 -75
rect 106 -87 115 -77
rect 73 -93 80 -87
rect 108 -93 115 -87
rect 117 -93 122 -73
rect 124 -80 129 -73
rect 167 -76 172 -73
rect 157 -79 162 -76
rect 124 -82 131 -80
rect 124 -84 127 -82
rect 129 -84 131 -82
rect 124 -86 131 -84
rect 135 -82 142 -79
rect 135 -84 137 -82
rect 139 -84 142 -82
rect 124 -93 129 -86
rect 135 -89 142 -84
rect 135 -91 137 -89
rect 139 -91 142 -89
rect 135 -93 142 -91
rect 144 -89 152 -79
rect 144 -91 147 -89
rect 149 -91 152 -89
rect 144 -93 152 -91
rect 154 -81 162 -79
rect 154 -83 157 -81
rect 159 -83 162 -81
rect 154 -86 162 -83
rect 164 -78 172 -76
rect 164 -80 167 -78
rect 169 -80 172 -78
rect 164 -86 172 -80
rect 174 -80 179 -73
rect 186 -76 192 -74
rect 186 -78 188 -76
rect 190 -78 192 -76
rect 186 -80 192 -78
rect 205 -76 211 -74
rect 205 -78 207 -76
rect 209 -78 211 -76
rect 205 -80 211 -78
rect 174 -82 181 -80
rect 174 -84 177 -82
rect 179 -84 181 -82
rect 174 -86 181 -84
rect 154 -93 159 -86
rect 186 -87 191 -80
rect 207 -84 211 -80
rect 207 -87 213 -84
rect 186 -93 193 -87
rect 195 -89 203 -87
rect 195 -91 198 -89
rect 200 -91 203 -89
rect 195 -93 203 -91
rect 205 -93 213 -87
rect 215 -87 220 -84
rect 215 -89 222 -87
rect 215 -91 218 -89
rect 220 -91 222 -89
rect 215 -93 222 -91
<< pdif >>
rect 9 131 14 143
rect 7 129 14 131
rect 7 127 9 129
rect 11 127 14 129
rect 7 122 14 127
rect 7 120 9 122
rect 11 120 14 122
rect 7 118 14 120
rect 16 141 25 143
rect 16 139 20 141
rect 22 139 25 141
rect 48 141 62 143
rect 48 140 55 141
rect 16 131 25 139
rect 32 131 37 140
rect 16 118 27 131
rect 29 122 37 131
rect 29 120 32 122
rect 34 120 37 122
rect 29 118 37 120
rect 32 115 37 118
rect 39 115 44 140
rect 46 139 55 140
rect 57 139 62 141
rect 46 134 62 139
rect 46 132 55 134
rect 57 132 62 134
rect 46 115 62 132
rect 64 133 72 143
rect 64 131 67 133
rect 69 131 72 133
rect 64 126 72 131
rect 64 124 67 126
rect 69 124 72 126
rect 64 115 72 124
rect 74 141 82 143
rect 74 139 77 141
rect 79 139 82 141
rect 74 134 82 139
rect 74 132 77 134
rect 79 132 82 134
rect 74 115 82 132
rect 84 128 89 143
rect 99 128 104 143
rect 84 126 91 128
rect 84 124 87 126
rect 89 124 91 126
rect 84 119 91 124
rect 84 117 87 119
rect 89 117 91 119
rect 84 115 91 117
rect 97 126 104 128
rect 97 124 99 126
rect 101 124 104 126
rect 97 119 104 124
rect 97 117 99 119
rect 101 117 104 119
rect 97 115 104 117
rect 106 141 114 143
rect 106 139 109 141
rect 111 139 114 141
rect 106 134 114 139
rect 106 132 109 134
rect 111 132 114 134
rect 106 115 114 132
rect 116 133 124 143
rect 116 131 119 133
rect 121 131 124 133
rect 116 126 124 131
rect 116 124 119 126
rect 121 124 124 126
rect 116 115 124 124
rect 126 141 140 143
rect 126 139 131 141
rect 133 140 140 141
rect 163 141 172 143
rect 133 139 142 140
rect 126 134 142 139
rect 126 132 131 134
rect 133 132 142 134
rect 126 115 142 132
rect 144 115 149 140
rect 151 131 156 140
rect 163 139 166 141
rect 168 139 172 141
rect 163 131 172 139
rect 151 122 159 131
rect 151 120 154 122
rect 156 120 159 122
rect 151 118 159 120
rect 161 118 172 131
rect 174 131 179 143
rect 188 136 193 143
rect 186 134 193 136
rect 186 132 188 134
rect 190 132 193 134
rect 174 129 181 131
rect 186 130 193 132
rect 174 127 177 129
rect 179 127 181 129
rect 174 122 181 127
rect 188 122 193 130
rect 195 122 200 143
rect 202 141 211 143
rect 202 139 207 141
rect 209 139 211 141
rect 202 133 211 139
rect 202 122 213 133
rect 174 120 177 122
rect 179 120 181 122
rect 174 118 181 120
rect 151 115 156 118
rect 205 115 213 122
rect 215 131 222 133
rect 215 129 218 131
rect 220 129 222 131
rect 215 124 222 129
rect 215 122 218 124
rect 220 122 222 124
rect 215 120 222 122
rect 215 115 220 120
rect 32 36 37 39
rect 7 34 14 36
rect 7 32 9 34
rect 11 32 14 34
rect 7 27 14 32
rect 7 25 9 27
rect 11 25 14 27
rect 7 23 14 25
rect 9 11 14 23
rect 16 23 27 36
rect 29 34 37 36
rect 29 32 32 34
rect 34 32 37 34
rect 29 23 37 32
rect 16 15 25 23
rect 16 13 20 15
rect 22 13 25 15
rect 32 14 37 23
rect 39 14 44 39
rect 46 22 62 39
rect 46 20 55 22
rect 57 20 62 22
rect 46 15 62 20
rect 46 14 55 15
rect 16 11 25 13
rect 48 13 55 14
rect 57 13 62 15
rect 48 11 62 13
rect 64 30 72 39
rect 64 28 67 30
rect 69 28 72 30
rect 64 23 72 28
rect 64 21 67 23
rect 69 21 72 23
rect 64 11 72 21
rect 74 22 82 39
rect 74 20 77 22
rect 79 20 82 22
rect 74 15 82 20
rect 74 13 77 15
rect 79 13 82 15
rect 74 11 82 13
rect 84 37 91 39
rect 84 35 87 37
rect 89 35 91 37
rect 84 30 91 35
rect 84 28 87 30
rect 89 28 91 30
rect 84 26 91 28
rect 97 37 104 39
rect 97 35 99 37
rect 101 35 104 37
rect 97 30 104 35
rect 97 28 99 30
rect 101 28 104 30
rect 97 26 104 28
rect 84 11 89 26
rect 99 11 104 26
rect 106 22 114 39
rect 106 20 109 22
rect 111 20 114 22
rect 106 15 114 20
rect 106 13 109 15
rect 111 13 114 15
rect 106 11 114 13
rect 116 30 124 39
rect 116 28 119 30
rect 121 28 124 30
rect 116 23 124 28
rect 116 21 119 23
rect 121 21 124 23
rect 116 11 124 21
rect 126 22 142 39
rect 126 20 131 22
rect 133 20 142 22
rect 126 15 142 20
rect 126 13 131 15
rect 133 14 142 15
rect 144 14 149 39
rect 151 36 156 39
rect 151 34 159 36
rect 151 32 154 34
rect 156 32 159 34
rect 151 23 159 32
rect 161 23 172 36
rect 151 14 156 23
rect 163 15 172 23
rect 133 13 140 14
rect 126 11 140 13
rect 163 13 166 15
rect 168 13 172 15
rect 163 11 172 13
rect 174 34 181 36
rect 174 32 177 34
rect 179 32 181 34
rect 205 32 213 39
rect 174 27 181 32
rect 174 25 177 27
rect 179 25 181 27
rect 174 23 181 25
rect 188 24 193 32
rect 174 11 179 23
rect 186 22 193 24
rect 186 20 188 22
rect 190 20 193 22
rect 186 18 193 20
rect 188 11 193 18
rect 195 11 200 32
rect 202 21 213 32
rect 215 34 220 39
rect 215 32 222 34
rect 215 30 218 32
rect 220 30 222 32
rect 215 25 222 30
rect 215 23 218 25
rect 220 23 222 25
rect 215 21 222 23
rect 202 15 211 21
rect 202 13 207 15
rect 209 13 211 15
rect 202 11 211 13
rect 9 -13 14 -1
rect 7 -15 14 -13
rect 7 -17 9 -15
rect 11 -17 14 -15
rect 7 -22 14 -17
rect 7 -24 9 -22
rect 11 -24 14 -22
rect 7 -26 14 -24
rect 16 -3 25 -1
rect 16 -5 20 -3
rect 22 -5 25 -3
rect 48 -3 62 -1
rect 48 -4 55 -3
rect 16 -13 25 -5
rect 32 -13 37 -4
rect 16 -26 27 -13
rect 29 -22 37 -13
rect 29 -24 32 -22
rect 34 -24 37 -22
rect 29 -26 37 -24
rect 32 -29 37 -26
rect 39 -29 44 -4
rect 46 -5 55 -4
rect 57 -5 62 -3
rect 46 -10 62 -5
rect 46 -12 55 -10
rect 57 -12 62 -10
rect 46 -29 62 -12
rect 64 -11 72 -1
rect 64 -13 67 -11
rect 69 -13 72 -11
rect 64 -18 72 -13
rect 64 -20 67 -18
rect 69 -20 72 -18
rect 64 -29 72 -20
rect 74 -3 82 -1
rect 74 -5 77 -3
rect 79 -5 82 -3
rect 74 -10 82 -5
rect 74 -12 77 -10
rect 79 -12 82 -10
rect 74 -29 82 -12
rect 84 -16 89 -1
rect 99 -16 104 -1
rect 84 -18 91 -16
rect 84 -20 87 -18
rect 89 -20 91 -18
rect 84 -25 91 -20
rect 84 -27 87 -25
rect 89 -27 91 -25
rect 84 -29 91 -27
rect 97 -18 104 -16
rect 97 -20 99 -18
rect 101 -20 104 -18
rect 97 -25 104 -20
rect 97 -27 99 -25
rect 101 -27 104 -25
rect 97 -29 104 -27
rect 106 -3 114 -1
rect 106 -5 109 -3
rect 111 -5 114 -3
rect 106 -10 114 -5
rect 106 -12 109 -10
rect 111 -12 114 -10
rect 106 -29 114 -12
rect 116 -11 124 -1
rect 116 -13 119 -11
rect 121 -13 124 -11
rect 116 -18 124 -13
rect 116 -20 119 -18
rect 121 -20 124 -18
rect 116 -29 124 -20
rect 126 -3 140 -1
rect 126 -5 131 -3
rect 133 -4 140 -3
rect 163 -3 172 -1
rect 133 -5 142 -4
rect 126 -10 142 -5
rect 126 -12 131 -10
rect 133 -12 142 -10
rect 126 -29 142 -12
rect 144 -29 149 -4
rect 151 -13 156 -4
rect 163 -5 166 -3
rect 168 -5 172 -3
rect 163 -13 172 -5
rect 151 -22 159 -13
rect 151 -24 154 -22
rect 156 -24 159 -22
rect 151 -26 159 -24
rect 161 -26 172 -13
rect 174 -13 179 -1
rect 188 -8 193 -1
rect 186 -10 193 -8
rect 186 -12 188 -10
rect 190 -12 193 -10
rect 174 -15 181 -13
rect 186 -14 193 -12
rect 174 -17 177 -15
rect 179 -17 181 -15
rect 174 -22 181 -17
rect 188 -22 193 -14
rect 195 -22 200 -1
rect 202 -3 211 -1
rect 202 -5 207 -3
rect 209 -5 211 -3
rect 202 -11 211 -5
rect 202 -22 213 -11
rect 174 -24 177 -22
rect 179 -24 181 -22
rect 174 -26 181 -24
rect 151 -29 156 -26
rect 205 -29 213 -22
rect 215 -13 222 -11
rect 215 -15 218 -13
rect 220 -15 222 -13
rect 215 -20 222 -15
rect 215 -22 218 -20
rect 220 -22 222 -20
rect 215 -24 222 -22
rect 215 -29 220 -24
rect 32 -108 37 -105
rect 7 -110 14 -108
rect 7 -112 9 -110
rect 11 -112 14 -110
rect 7 -117 14 -112
rect 7 -119 9 -117
rect 11 -119 14 -117
rect 7 -121 14 -119
rect 9 -133 14 -121
rect 16 -121 27 -108
rect 29 -110 37 -108
rect 29 -112 32 -110
rect 34 -112 37 -110
rect 29 -121 37 -112
rect 16 -129 25 -121
rect 16 -131 20 -129
rect 22 -131 25 -129
rect 32 -130 37 -121
rect 39 -130 44 -105
rect 46 -122 62 -105
rect 46 -124 55 -122
rect 57 -124 62 -122
rect 46 -129 62 -124
rect 46 -130 55 -129
rect 16 -133 25 -131
rect 48 -131 55 -130
rect 57 -131 62 -129
rect 48 -133 62 -131
rect 64 -114 72 -105
rect 64 -116 67 -114
rect 69 -116 72 -114
rect 64 -121 72 -116
rect 64 -123 67 -121
rect 69 -123 72 -121
rect 64 -133 72 -123
rect 74 -122 82 -105
rect 74 -124 77 -122
rect 79 -124 82 -122
rect 74 -129 82 -124
rect 74 -131 77 -129
rect 79 -131 82 -129
rect 74 -133 82 -131
rect 84 -107 91 -105
rect 84 -109 87 -107
rect 89 -109 91 -107
rect 84 -114 91 -109
rect 84 -116 87 -114
rect 89 -116 91 -114
rect 84 -118 91 -116
rect 97 -107 104 -105
rect 97 -109 99 -107
rect 101 -109 104 -107
rect 97 -114 104 -109
rect 97 -116 99 -114
rect 101 -116 104 -114
rect 97 -118 104 -116
rect 84 -133 89 -118
rect 99 -133 104 -118
rect 106 -122 114 -105
rect 106 -124 109 -122
rect 111 -124 114 -122
rect 106 -129 114 -124
rect 106 -131 109 -129
rect 111 -131 114 -129
rect 106 -133 114 -131
rect 116 -114 124 -105
rect 116 -116 119 -114
rect 121 -116 124 -114
rect 116 -121 124 -116
rect 116 -123 119 -121
rect 121 -123 124 -121
rect 116 -133 124 -123
rect 126 -122 142 -105
rect 126 -124 131 -122
rect 133 -124 142 -122
rect 126 -129 142 -124
rect 126 -131 131 -129
rect 133 -130 142 -129
rect 144 -130 149 -105
rect 151 -108 156 -105
rect 151 -110 159 -108
rect 151 -112 154 -110
rect 156 -112 159 -110
rect 151 -121 159 -112
rect 161 -121 172 -108
rect 151 -130 156 -121
rect 163 -129 172 -121
rect 133 -131 140 -130
rect 126 -133 140 -131
rect 163 -131 166 -129
rect 168 -131 172 -129
rect 163 -133 172 -131
rect 174 -110 181 -108
rect 174 -112 177 -110
rect 179 -112 181 -110
rect 205 -112 213 -105
rect 174 -117 181 -112
rect 174 -119 177 -117
rect 179 -119 181 -117
rect 174 -121 181 -119
rect 188 -120 193 -112
rect 174 -133 179 -121
rect 186 -122 193 -120
rect 186 -124 188 -122
rect 190 -124 193 -122
rect 186 -126 193 -124
rect 188 -133 193 -126
rect 195 -133 200 -112
rect 202 -123 213 -112
rect 215 -110 220 -105
rect 215 -112 222 -110
rect 215 -114 218 -112
rect 220 -114 222 -112
rect 215 -119 222 -114
rect 215 -121 218 -119
rect 220 -121 222 -119
rect 215 -123 222 -121
rect 202 -129 211 -123
rect 202 -131 207 -129
rect 209 -131 211 -129
rect 202 -133 211 -131
<< alu1 >>
rect 3 144 225 149
rect 3 142 217 144
rect 219 142 225 144
rect 3 141 225 142
rect 218 135 222 136
rect 209 131 222 135
rect 7 129 12 131
rect 7 127 9 129
rect 11 127 12 129
rect 7 122 12 127
rect 7 120 9 122
rect 11 120 12 122
rect 7 118 12 120
rect 7 102 11 118
rect 38 115 76 119
rect 38 112 43 115
rect 35 110 43 112
rect 35 108 36 110
rect 38 108 43 110
rect 35 106 43 108
rect 53 110 68 111
rect 53 108 55 110
rect 57 108 62 110
rect 64 108 68 110
rect 53 107 68 108
rect 7 100 8 102
rect 10 100 11 102
rect 7 96 11 100
rect 7 94 12 96
rect 55 98 59 107
rect 86 126 92 128
rect 86 124 87 126
rect 89 124 92 126
rect 86 119 92 124
rect 86 117 87 119
rect 89 117 92 119
rect 86 115 92 117
rect 88 110 92 115
rect 88 108 89 110
rect 91 108 92 110
rect 88 95 92 108
rect 7 92 9 94
rect 11 92 12 94
rect 7 90 12 92
rect 86 94 92 95
rect 86 92 87 94
rect 89 92 92 94
rect 86 91 92 92
rect 96 126 102 128
rect 176 129 181 131
rect 176 127 177 129
rect 179 127 181 129
rect 96 124 99 126
rect 101 124 102 126
rect 96 123 102 124
rect 96 121 99 123
rect 101 121 102 123
rect 96 119 102 121
rect 96 117 99 119
rect 101 117 102 119
rect 96 115 102 117
rect 96 95 100 115
rect 112 115 150 119
rect 145 112 150 115
rect 120 110 135 111
rect 120 108 124 110
rect 126 108 131 110
rect 133 108 135 110
rect 120 107 135 108
rect 145 110 153 112
rect 145 108 150 110
rect 152 108 153 110
rect 129 102 133 107
rect 145 106 153 108
rect 176 122 181 127
rect 176 120 177 122
rect 179 120 181 122
rect 176 118 181 120
rect 129 100 130 102
rect 132 100 133 102
rect 129 98 133 100
rect 96 94 102 95
rect 96 92 99 94
rect 101 92 102 94
rect 96 91 102 92
rect 177 96 181 118
rect 186 123 190 128
rect 186 121 187 123
rect 189 121 190 123
rect 186 119 190 121
rect 186 117 207 119
rect 186 115 191 117
rect 193 115 207 117
rect 186 110 207 111
rect 186 108 187 110
rect 189 108 201 110
rect 203 108 207 110
rect 186 107 207 108
rect 220 129 222 131
rect 218 124 222 129
rect 220 122 222 124
rect 186 98 190 107
rect 218 106 222 122
rect 218 104 219 106
rect 221 104 222 106
rect 218 103 222 104
rect 217 101 222 103
rect 217 99 218 101
rect 220 99 222 101
rect 217 97 222 99
rect 176 94 181 96
rect 176 92 177 94
rect 179 92 181 94
rect 176 90 181 92
rect 3 84 225 85
rect 3 82 217 84
rect 219 82 225 84
rect 3 72 225 82
rect 3 70 217 72
rect 219 70 225 72
rect 3 69 225 70
rect 7 62 12 64
rect 7 60 9 62
rect 11 60 12 62
rect 7 58 12 60
rect 7 54 11 58
rect 7 52 8 54
rect 10 52 11 54
rect 7 36 11 52
rect 86 62 92 63
rect 86 60 87 62
rect 89 60 92 62
rect 86 59 92 60
rect 7 34 12 36
rect 7 32 9 34
rect 11 32 12 34
rect 7 27 12 32
rect 35 46 43 48
rect 55 47 59 56
rect 35 44 36 46
rect 38 44 43 46
rect 35 42 43 44
rect 53 46 68 47
rect 53 44 55 46
rect 57 44 62 46
rect 64 44 68 46
rect 53 43 68 44
rect 38 39 43 42
rect 88 46 92 59
rect 88 44 89 46
rect 91 44 92 46
rect 38 35 76 39
rect 88 39 92 44
rect 86 37 92 39
rect 86 35 87 37
rect 89 35 92 37
rect 86 30 92 35
rect 86 28 87 30
rect 89 28 92 30
rect 7 25 9 27
rect 11 25 12 27
rect 7 23 12 25
rect 86 26 92 28
rect 96 62 102 63
rect 96 60 99 62
rect 101 60 102 62
rect 96 59 102 60
rect 176 62 181 64
rect 176 60 177 62
rect 179 60 181 62
rect 96 39 100 59
rect 129 54 133 56
rect 129 52 130 54
rect 132 52 133 54
rect 96 37 102 39
rect 96 35 99 37
rect 101 35 102 37
rect 96 33 102 35
rect 96 31 99 33
rect 101 31 102 33
rect 96 30 102 31
rect 96 28 99 30
rect 101 28 102 30
rect 96 26 102 28
rect 129 47 133 52
rect 176 58 181 60
rect 120 46 135 47
rect 120 44 124 46
rect 126 44 131 46
rect 133 44 135 46
rect 120 43 135 44
rect 145 46 153 48
rect 145 44 150 46
rect 152 44 153 46
rect 145 42 153 44
rect 145 41 150 42
rect 145 39 147 41
rect 149 39 150 41
rect 112 35 150 39
rect 177 36 181 58
rect 186 52 190 56
rect 186 50 187 52
rect 189 50 190 52
rect 186 47 190 50
rect 186 46 207 47
rect 186 44 201 46
rect 203 44 207 46
rect 186 43 207 44
rect 217 55 222 57
rect 217 53 218 55
rect 220 53 222 55
rect 217 51 222 53
rect 176 34 181 36
rect 176 32 177 34
rect 179 32 181 34
rect 176 27 181 32
rect 176 25 177 27
rect 179 25 181 27
rect 186 37 191 39
rect 193 37 207 39
rect 186 35 207 37
rect 186 33 190 35
rect 186 31 187 33
rect 189 31 190 33
rect 186 26 190 31
rect 176 23 181 25
rect 218 32 222 51
rect 220 30 222 32
rect 218 25 222 30
rect 220 23 222 25
rect 209 22 222 23
rect 209 20 211 22
rect 213 20 222 22
rect 209 19 222 20
rect 218 18 222 19
rect 3 12 225 13
rect 3 10 217 12
rect 219 10 225 12
rect 3 0 225 10
rect 3 -2 217 0
rect 219 -2 225 0
rect 3 -3 225 -2
rect 218 -9 222 -8
rect 209 -13 222 -9
rect 7 -15 12 -13
rect 7 -17 9 -15
rect 11 -17 12 -15
rect 7 -22 12 -17
rect 7 -24 9 -22
rect 11 -24 12 -22
rect 7 -26 12 -24
rect 7 -42 11 -26
rect 38 -29 76 -25
rect 38 -32 43 -29
rect 35 -34 43 -32
rect 35 -36 36 -34
rect 38 -36 43 -34
rect 35 -38 43 -36
rect 53 -34 68 -33
rect 53 -36 55 -34
rect 57 -36 62 -34
rect 64 -36 68 -34
rect 53 -37 68 -36
rect 7 -44 8 -42
rect 10 -44 11 -42
rect 7 -48 11 -44
rect 7 -50 12 -48
rect 55 -46 59 -37
rect 86 -18 92 -16
rect 86 -20 87 -18
rect 89 -20 92 -18
rect 86 -25 92 -20
rect 86 -27 87 -25
rect 89 -27 92 -25
rect 86 -29 92 -27
rect 88 -34 92 -29
rect 88 -36 89 -34
rect 91 -36 92 -34
rect 88 -49 92 -36
rect 7 -52 9 -50
rect 11 -52 12 -50
rect 7 -54 12 -52
rect 86 -50 92 -49
rect 86 -52 87 -50
rect 89 -52 92 -50
rect 86 -53 92 -52
rect 96 -18 102 -16
rect 176 -15 181 -13
rect 176 -17 177 -15
rect 179 -17 181 -15
rect 96 -20 99 -18
rect 101 -20 102 -18
rect 96 -21 102 -20
rect 96 -23 99 -21
rect 101 -23 102 -21
rect 96 -25 102 -23
rect 96 -27 99 -25
rect 101 -27 102 -25
rect 96 -29 102 -27
rect 96 -49 100 -29
rect 112 -26 150 -25
rect 112 -28 147 -26
rect 149 -28 150 -26
rect 112 -29 150 -28
rect 145 -32 150 -29
rect 120 -34 135 -33
rect 120 -36 124 -34
rect 126 -36 131 -34
rect 133 -36 135 -34
rect 120 -37 135 -36
rect 145 -34 153 -32
rect 145 -36 150 -34
rect 152 -36 153 -34
rect 129 -42 133 -37
rect 145 -38 153 -36
rect 176 -22 181 -17
rect 176 -24 177 -22
rect 179 -24 181 -22
rect 176 -26 181 -24
rect 129 -44 130 -42
rect 132 -44 133 -42
rect 129 -46 133 -44
rect 96 -50 102 -49
rect 96 -52 99 -50
rect 101 -52 102 -50
rect 96 -53 102 -52
rect 177 -48 181 -26
rect 186 -17 190 -16
rect 186 -19 187 -17
rect 189 -19 190 -17
rect 186 -25 190 -19
rect 186 -27 207 -25
rect 186 -29 191 -27
rect 193 -29 207 -27
rect 186 -34 207 -33
rect 186 -36 187 -34
rect 189 -36 201 -34
rect 203 -36 207 -34
rect 186 -37 207 -36
rect 220 -15 222 -13
rect 218 -20 222 -15
rect 220 -22 222 -20
rect 186 -46 190 -37
rect 218 -38 222 -22
rect 218 -40 219 -38
rect 221 -40 222 -38
rect 218 -41 222 -40
rect 217 -43 222 -41
rect 217 -45 218 -43
rect 220 -45 222 -43
rect 217 -47 222 -45
rect 176 -50 181 -48
rect 176 -52 177 -50
rect 179 -52 181 -50
rect 176 -54 181 -52
rect 3 -60 225 -59
rect 3 -62 217 -60
rect 219 -62 225 -60
rect 3 -72 225 -62
rect 3 -74 217 -72
rect 219 -74 225 -72
rect 3 -75 225 -74
rect 7 -82 12 -80
rect 7 -84 9 -82
rect 11 -84 12 -82
rect 7 -86 12 -84
rect 7 -90 11 -86
rect 7 -92 8 -90
rect 10 -92 11 -90
rect 7 -108 11 -92
rect 86 -82 92 -81
rect 86 -84 87 -82
rect 89 -84 92 -82
rect 86 -85 92 -84
rect 7 -110 12 -108
rect 7 -112 9 -110
rect 11 -112 12 -110
rect 7 -117 12 -112
rect 35 -98 43 -96
rect 55 -97 59 -88
rect 35 -100 36 -98
rect 38 -100 43 -98
rect 35 -102 43 -100
rect 53 -98 68 -97
rect 53 -100 55 -98
rect 57 -100 62 -98
rect 64 -100 68 -98
rect 53 -101 68 -100
rect 38 -105 43 -102
rect 88 -98 92 -85
rect 88 -100 89 -98
rect 91 -100 92 -98
rect 38 -109 76 -105
rect 88 -105 92 -100
rect 86 -107 92 -105
rect 86 -109 87 -107
rect 89 -109 92 -107
rect 86 -114 92 -109
rect 86 -116 87 -114
rect 89 -116 92 -114
rect 7 -119 9 -117
rect 11 -119 12 -117
rect 7 -121 12 -119
rect 86 -118 92 -116
rect 96 -82 102 -81
rect 96 -84 99 -82
rect 101 -84 102 -82
rect 96 -85 102 -84
rect 176 -82 181 -80
rect 176 -84 177 -82
rect 179 -84 181 -82
rect 96 -105 100 -85
rect 129 -90 133 -88
rect 129 -92 130 -90
rect 132 -92 133 -90
rect 96 -107 102 -105
rect 96 -109 99 -107
rect 101 -109 102 -107
rect 96 -111 102 -109
rect 96 -113 99 -111
rect 101 -113 102 -111
rect 96 -114 102 -113
rect 96 -116 99 -114
rect 101 -116 102 -114
rect 96 -118 102 -116
rect 129 -97 133 -92
rect 176 -86 181 -84
rect 120 -98 135 -97
rect 120 -100 124 -98
rect 126 -100 131 -98
rect 133 -100 135 -98
rect 120 -101 135 -100
rect 145 -98 153 -96
rect 145 -100 150 -98
rect 152 -100 153 -98
rect 145 -102 153 -100
rect 145 -103 150 -102
rect 145 -105 147 -103
rect 149 -105 150 -103
rect 112 -109 150 -105
rect 177 -108 181 -86
rect 186 -92 190 -88
rect 186 -94 187 -92
rect 189 -94 190 -92
rect 186 -97 190 -94
rect 186 -98 207 -97
rect 186 -100 201 -98
rect 203 -100 207 -98
rect 186 -101 207 -100
rect 217 -89 222 -87
rect 217 -91 218 -89
rect 220 -91 222 -89
rect 217 -93 222 -91
rect 176 -110 181 -108
rect 176 -112 177 -110
rect 179 -112 181 -110
rect 176 -117 181 -112
rect 176 -119 177 -117
rect 179 -119 181 -117
rect 186 -107 191 -105
rect 193 -107 207 -105
rect 186 -109 207 -107
rect 186 -111 190 -109
rect 186 -113 187 -111
rect 189 -113 190 -111
rect 186 -118 190 -113
rect 176 -121 181 -119
rect 218 -112 222 -93
rect 220 -114 222 -112
rect 218 -119 222 -114
rect 220 -121 222 -119
rect 209 -125 222 -121
rect 218 -126 222 -125
rect 3 -132 225 -131
rect 3 -134 217 -132
rect 219 -134 225 -132
rect 3 -139 225 -134
<< alu2 >>
rect 98 123 190 124
rect 98 121 99 123
rect 101 121 187 123
rect 189 121 190 123
rect 98 120 190 121
rect 88 110 191 111
rect 88 108 89 110
rect 91 108 187 110
rect 189 108 191 110
rect 88 107 191 108
rect 218 106 226 107
rect 218 104 219 106
rect 221 104 223 106
rect 225 104 226 106
rect 218 103 226 104
rect 7 102 133 103
rect 7 100 8 102
rect 10 100 130 102
rect 132 100 133 102
rect 7 99 133 100
rect 7 54 133 55
rect 7 52 8 54
rect 10 52 130 54
rect 132 52 133 54
rect 7 51 133 52
rect 137 52 190 53
rect 137 50 187 52
rect 189 50 190 52
rect 137 49 190 50
rect 137 47 141 49
rect 88 46 141 47
rect 88 44 89 46
rect 91 44 141 46
rect 88 43 141 44
rect 146 41 226 42
rect 146 39 147 41
rect 149 39 223 41
rect 225 39 226 41
rect 146 38 226 39
rect 98 33 190 34
rect 98 31 99 33
rect 101 31 187 33
rect 189 31 190 33
rect 98 30 190 31
rect 210 22 214 23
rect 210 20 211 22
rect 213 20 214 22
rect 138 -17 190 -16
rect 138 -19 187 -17
rect 189 -19 190 -17
rect 138 -20 190 -19
rect 98 -21 142 -20
rect 98 -23 99 -21
rect 101 -23 142 -21
rect 98 -24 142 -23
rect 210 -25 214 20
rect 146 -26 214 -25
rect 146 -28 147 -26
rect 149 -28 214 -26
rect 146 -29 214 -28
rect 88 -34 191 -33
rect 88 -36 89 -34
rect 91 -36 187 -34
rect 189 -36 191 -34
rect 88 -37 191 -36
rect 218 -38 226 -37
rect 218 -40 219 -38
rect 221 -40 223 -38
rect 225 -40 226 -38
rect 218 -41 226 -40
rect 7 -42 133 -41
rect 7 -44 8 -42
rect 10 -44 130 -42
rect 132 -44 133 -42
rect 7 -45 133 -44
rect 7 -90 133 -89
rect 7 -92 8 -90
rect 10 -92 130 -90
rect 132 -92 133 -90
rect 7 -93 133 -92
rect 137 -92 190 -91
rect 137 -94 187 -92
rect 189 -94 190 -92
rect 137 -95 190 -94
rect 137 -97 141 -95
rect 88 -98 141 -97
rect 88 -100 89 -98
rect 91 -100 141 -98
rect 88 -101 141 -100
rect 146 -103 226 -102
rect 146 -105 147 -103
rect 149 -105 223 -103
rect 225 -105 226 -103
rect 146 -106 226 -105
rect 98 -111 190 -110
rect 98 -113 99 -111
rect 101 -113 187 -111
rect 189 -113 190 -111
rect 98 -114 190 -113
<< alu3 >>
rect 222 106 226 107
rect 222 104 223 106
rect 225 104 226 106
rect 222 41 226 104
rect 222 39 223 41
rect 225 39 226 41
rect 222 38 226 39
rect 222 -38 226 -37
rect 222 -40 223 -38
rect 225 -40 226 -38
rect 222 -103 226 -40
rect 222 -105 223 -103
rect 225 -105 226 -103
rect 222 -106 226 -105
<< ptie >>
rect 215 84 221 86
rect 215 82 217 84
rect 219 82 221 84
rect 215 80 221 82
rect 215 72 221 74
rect 215 70 217 72
rect 219 70 221 72
rect 215 68 221 70
rect 215 -60 221 -58
rect 215 -62 217 -60
rect 219 -62 221 -60
rect 215 -64 221 -62
rect 215 -72 221 -70
rect 215 -74 217 -72
rect 219 -74 221 -72
rect 215 -76 221 -74
<< ntie >>
rect 215 144 221 146
rect 215 142 217 144
rect 219 142 221 144
rect 215 140 221 142
rect 215 12 221 14
rect 215 10 217 12
rect 219 10 221 12
rect 215 8 221 10
rect 215 0 221 2
rect 215 -2 217 0
rect 219 -2 221 0
rect 215 -4 221 -2
rect 215 -132 221 -130
rect 215 -134 217 -132
rect 219 -134 221 -132
rect 215 -136 221 -134
<< nmos >>
rect 14 83 16 96
rect 24 86 26 96
rect 34 89 36 103
rect 44 89 46 103
rect 64 83 66 103
rect 71 83 73 103
rect 82 83 84 97
rect 104 83 106 97
rect 115 83 117 103
rect 122 83 124 103
rect 142 89 144 103
rect 152 89 154 103
rect 193 97 195 103
rect 203 97 205 103
rect 162 86 164 96
rect 172 83 174 96
rect 213 94 215 103
rect 14 58 16 71
rect 24 58 26 68
rect 34 51 36 65
rect 44 51 46 65
rect 64 51 66 71
rect 71 51 73 71
rect 82 57 84 71
rect 104 57 106 71
rect 115 51 117 71
rect 122 51 124 71
rect 142 51 144 65
rect 152 51 154 65
rect 162 58 164 68
rect 172 58 174 71
rect 193 51 195 57
rect 203 51 205 57
rect 213 51 215 60
rect 14 -61 16 -48
rect 24 -58 26 -48
rect 34 -55 36 -41
rect 44 -55 46 -41
rect 64 -61 66 -41
rect 71 -61 73 -41
rect 82 -61 84 -47
rect 104 -61 106 -47
rect 115 -61 117 -41
rect 122 -61 124 -41
rect 142 -55 144 -41
rect 152 -55 154 -41
rect 193 -47 195 -41
rect 203 -47 205 -41
rect 162 -58 164 -48
rect 172 -61 174 -48
rect 213 -50 215 -41
rect 14 -86 16 -73
rect 24 -86 26 -76
rect 34 -93 36 -79
rect 44 -93 46 -79
rect 64 -93 66 -73
rect 71 -93 73 -73
rect 82 -87 84 -73
rect 104 -87 106 -73
rect 115 -93 117 -73
rect 122 -93 124 -73
rect 142 -93 144 -79
rect 152 -93 154 -79
rect 162 -86 164 -76
rect 172 -86 174 -73
rect 193 -93 195 -87
rect 203 -93 205 -87
rect 213 -93 215 -84
<< pmos >>
rect 14 118 16 143
rect 27 118 29 131
rect 37 115 39 140
rect 44 115 46 140
rect 62 115 64 143
rect 72 115 74 143
rect 82 115 84 143
rect 104 115 106 143
rect 114 115 116 143
rect 124 115 126 143
rect 142 115 144 140
rect 149 115 151 140
rect 159 118 161 131
rect 172 118 174 143
rect 193 122 195 143
rect 200 122 202 143
rect 213 115 215 133
rect 14 11 16 36
rect 27 23 29 36
rect 37 14 39 39
rect 44 14 46 39
rect 62 11 64 39
rect 72 11 74 39
rect 82 11 84 39
rect 104 11 106 39
rect 114 11 116 39
rect 124 11 126 39
rect 142 14 144 39
rect 149 14 151 39
rect 159 23 161 36
rect 172 11 174 36
rect 193 11 195 32
rect 200 11 202 32
rect 213 21 215 39
rect 14 -26 16 -1
rect 27 -26 29 -13
rect 37 -29 39 -4
rect 44 -29 46 -4
rect 62 -29 64 -1
rect 72 -29 74 -1
rect 82 -29 84 -1
rect 104 -29 106 -1
rect 114 -29 116 -1
rect 124 -29 126 -1
rect 142 -29 144 -4
rect 149 -29 151 -4
rect 159 -26 161 -13
rect 172 -26 174 -1
rect 193 -22 195 -1
rect 200 -22 202 -1
rect 213 -29 215 -11
rect 14 -133 16 -108
rect 27 -121 29 -108
rect 37 -130 39 -105
rect 44 -130 46 -105
rect 62 -133 64 -105
rect 72 -133 74 -105
rect 82 -133 84 -105
rect 104 -133 106 -105
rect 114 -133 116 -105
rect 124 -133 126 -105
rect 142 -130 144 -105
rect 149 -130 151 -105
rect 159 -121 161 -108
rect 172 -133 174 -108
rect 193 -133 195 -112
rect 200 -133 202 -112
rect 213 -123 215 -105
<< polyct0 >>
rect 22 111 24 113
rect 16 101 18 103
rect 72 108 74 110
rect 82 108 84 110
rect 104 108 106 110
rect 114 108 116 110
rect 164 111 166 113
rect 211 108 213 110
rect 170 101 172 103
rect 16 51 18 53
rect 22 41 24 43
rect 72 44 74 46
rect 82 44 84 46
rect 104 44 106 46
rect 114 44 116 46
rect 170 51 172 53
rect 164 41 166 43
rect 211 44 213 46
rect 22 -33 24 -31
rect 16 -43 18 -41
rect 72 -36 74 -34
rect 82 -36 84 -34
rect 104 -36 106 -34
rect 114 -36 116 -34
rect 164 -33 166 -31
rect 211 -36 213 -34
rect 170 -43 172 -41
rect 16 -93 18 -91
rect 22 -103 24 -101
rect 72 -100 74 -98
rect 82 -100 84 -98
rect 104 -100 106 -98
rect 114 -100 116 -98
rect 170 -93 172 -91
rect 164 -103 166 -101
rect 211 -100 213 -98
<< polyct1 >>
rect 36 108 38 110
rect 55 108 57 110
rect 62 108 64 110
rect 124 108 126 110
rect 131 108 133 110
rect 150 108 152 110
rect 191 115 193 117
rect 201 108 203 110
rect 36 44 38 46
rect 55 44 57 46
rect 62 44 64 46
rect 124 44 126 46
rect 131 44 133 46
rect 150 44 152 46
rect 201 44 203 46
rect 191 37 193 39
rect 36 -36 38 -34
rect 55 -36 57 -34
rect 62 -36 64 -34
rect 124 -36 126 -34
rect 131 -36 133 -34
rect 150 -36 152 -34
rect 191 -29 193 -27
rect 201 -36 203 -34
rect 36 -100 38 -98
rect 55 -100 57 -98
rect 62 -100 64 -98
rect 124 -100 126 -98
rect 131 -100 133 -98
rect 150 -100 152 -98
rect 201 -100 203 -98
rect 191 -107 193 -105
<< ndifct0 >>
rect 19 88 21 90
rect 29 91 31 93
rect 39 99 41 101
rect 49 99 51 101
rect 49 92 51 94
rect 59 92 61 94
rect 76 85 78 87
rect 110 85 112 87
rect 137 99 139 101
rect 127 92 129 94
rect 137 92 139 94
rect 147 99 149 101
rect 198 99 200 101
rect 157 91 159 93
rect 167 88 169 90
rect 188 86 190 88
rect 207 86 209 88
rect 19 64 21 66
rect 29 61 31 63
rect 39 53 41 55
rect 49 60 51 62
rect 59 60 61 62
rect 49 53 51 55
rect 76 67 78 69
rect 110 67 112 69
rect 127 60 129 62
rect 137 60 139 62
rect 137 53 139 55
rect 147 53 149 55
rect 157 61 159 63
rect 167 64 169 66
rect 188 66 190 68
rect 207 66 209 68
rect 198 53 200 55
rect 19 -56 21 -54
rect 29 -53 31 -51
rect 39 -45 41 -43
rect 49 -45 51 -43
rect 49 -52 51 -50
rect 59 -52 61 -50
rect 76 -59 78 -57
rect 110 -59 112 -57
rect 137 -45 139 -43
rect 127 -52 129 -50
rect 137 -52 139 -50
rect 147 -45 149 -43
rect 198 -45 200 -43
rect 157 -53 159 -51
rect 167 -56 169 -54
rect 188 -58 190 -56
rect 207 -58 209 -56
rect 19 -80 21 -78
rect 29 -83 31 -81
rect 39 -91 41 -89
rect 49 -84 51 -82
rect 59 -84 61 -82
rect 49 -91 51 -89
rect 76 -77 78 -75
rect 110 -77 112 -75
rect 127 -84 129 -82
rect 137 -84 139 -82
rect 137 -91 139 -89
rect 147 -91 149 -89
rect 157 -83 159 -81
rect 167 -80 169 -78
rect 188 -78 190 -76
rect 207 -78 209 -76
rect 198 -91 200 -89
<< ndifct1 >>
rect 9 92 11 94
rect 87 92 89 94
rect 99 92 101 94
rect 177 92 179 94
rect 218 99 220 101
rect 9 60 11 62
rect 87 60 89 62
rect 99 60 101 62
rect 177 60 179 62
rect 218 53 220 55
rect 9 -52 11 -50
rect 87 -52 89 -50
rect 99 -52 101 -50
rect 177 -52 179 -50
rect 218 -45 220 -43
rect 9 -84 11 -82
rect 87 -84 89 -82
rect 99 -84 101 -82
rect 177 -84 179 -82
rect 218 -91 220 -89
<< ntiect1 >>
rect 217 142 219 144
rect 217 10 219 12
rect 217 -2 219 0
rect 217 -134 219 -132
<< ptiect1 >>
rect 217 82 219 84
rect 217 70 219 72
rect 217 -62 219 -60
rect 217 -74 219 -72
<< pdifct0 >>
rect 20 139 22 141
rect 32 120 34 122
rect 55 139 57 141
rect 55 132 57 134
rect 67 131 69 133
rect 67 124 69 126
rect 77 139 79 141
rect 77 132 79 134
rect 109 139 111 141
rect 109 132 111 134
rect 119 131 121 133
rect 119 124 121 126
rect 131 139 133 141
rect 131 132 133 134
rect 166 139 168 141
rect 154 120 156 122
rect 188 132 190 134
rect 207 139 209 141
rect 32 32 34 34
rect 20 13 22 15
rect 55 20 57 22
rect 55 13 57 15
rect 67 28 69 30
rect 67 21 69 23
rect 77 20 79 22
rect 77 13 79 15
rect 109 20 111 22
rect 109 13 111 15
rect 119 28 121 30
rect 119 21 121 23
rect 131 20 133 22
rect 131 13 133 15
rect 154 32 156 34
rect 166 13 168 15
rect 188 20 190 22
rect 207 13 209 15
rect 20 -5 22 -3
rect 32 -24 34 -22
rect 55 -5 57 -3
rect 55 -12 57 -10
rect 67 -13 69 -11
rect 67 -20 69 -18
rect 77 -5 79 -3
rect 77 -12 79 -10
rect 109 -5 111 -3
rect 109 -12 111 -10
rect 119 -13 121 -11
rect 119 -20 121 -18
rect 131 -5 133 -3
rect 131 -12 133 -10
rect 166 -5 168 -3
rect 154 -24 156 -22
rect 188 -12 190 -10
rect 207 -5 209 -3
rect 32 -112 34 -110
rect 20 -131 22 -129
rect 55 -124 57 -122
rect 55 -131 57 -129
rect 67 -116 69 -114
rect 67 -123 69 -121
rect 77 -124 79 -122
rect 77 -131 79 -129
rect 109 -124 111 -122
rect 109 -131 111 -129
rect 119 -116 121 -114
rect 119 -123 121 -121
rect 131 -124 133 -122
rect 131 -131 133 -129
rect 154 -112 156 -110
rect 166 -131 168 -129
rect 188 -124 190 -122
rect 207 -131 209 -129
<< pdifct1 >>
rect 9 127 11 129
rect 9 120 11 122
rect 87 124 89 126
rect 87 117 89 119
rect 99 124 101 126
rect 99 117 101 119
rect 177 127 179 129
rect 177 120 179 122
rect 218 129 220 131
rect 218 122 220 124
rect 9 32 11 34
rect 9 25 11 27
rect 87 35 89 37
rect 87 28 89 30
rect 99 35 101 37
rect 99 28 101 30
rect 177 32 179 34
rect 177 25 179 27
rect 218 30 220 32
rect 218 23 220 25
rect 9 -17 11 -15
rect 9 -24 11 -22
rect 87 -20 89 -18
rect 87 -27 89 -25
rect 99 -20 101 -18
rect 99 -27 101 -25
rect 177 -17 179 -15
rect 177 -24 179 -22
rect 218 -15 220 -13
rect 218 -22 220 -20
rect 9 -112 11 -110
rect 9 -119 11 -117
rect 87 -109 89 -107
rect 87 -116 89 -114
rect 99 -109 101 -107
rect 99 -116 101 -114
rect 177 -112 179 -110
rect 177 -119 179 -117
rect 218 -114 220 -112
rect 218 -121 220 -119
<< alu0 >>
rect 18 139 20 141
rect 22 139 24 141
rect 18 138 24 139
rect 53 139 55 141
rect 57 139 59 141
rect 53 134 59 139
rect 75 139 77 141
rect 79 139 81 141
rect 53 132 55 134
rect 57 132 59 134
rect 53 131 59 132
rect 66 133 70 135
rect 66 131 67 133
rect 69 131 70 133
rect 75 134 81 139
rect 75 132 77 134
rect 79 132 81 134
rect 75 131 81 132
rect 107 139 109 141
rect 111 139 113 141
rect 107 134 113 139
rect 129 139 131 141
rect 133 139 135 141
rect 107 132 109 134
rect 111 132 113 134
rect 107 131 113 132
rect 118 133 122 135
rect 118 131 119 133
rect 121 131 122 133
rect 129 134 135 139
rect 164 139 166 141
rect 168 139 170 141
rect 164 138 170 139
rect 205 139 207 141
rect 209 139 211 141
rect 205 138 211 139
rect 129 132 131 134
rect 133 132 135 134
rect 129 131 135 132
rect 186 134 203 135
rect 186 132 188 134
rect 190 132 203 134
rect 186 131 203 132
rect 23 127 47 131
rect 66 127 70 131
rect 21 123 27 127
rect 43 126 83 127
rect 43 124 67 126
rect 69 124 83 126
rect 21 113 25 123
rect 31 122 35 124
rect 43 123 83 124
rect 31 120 32 122
rect 34 120 35 122
rect 31 119 35 120
rect 21 111 22 113
rect 24 111 25 113
rect 21 109 25 111
rect 28 115 35 119
rect 28 104 32 115
rect 71 110 75 115
rect 71 108 72 110
rect 74 108 75 110
rect 14 103 32 104
rect 14 101 16 103
rect 18 102 32 103
rect 18 101 43 102
rect 14 100 39 101
rect 28 99 39 100
rect 41 99 43 101
rect 28 98 43 99
rect 48 101 52 103
rect 48 99 49 101
rect 51 99 52 101
rect 48 94 52 99
rect 71 106 75 108
rect 79 112 83 123
rect 79 110 85 112
rect 79 108 82 110
rect 84 108 85 110
rect 79 106 85 108
rect 79 103 83 106
rect 63 99 83 103
rect 63 95 67 99
rect 27 93 49 94
rect 18 90 22 92
rect 27 91 29 93
rect 31 92 49 93
rect 51 92 52 94
rect 31 91 52 92
rect 57 94 67 95
rect 57 92 59 94
rect 61 92 67 94
rect 57 91 67 92
rect 118 127 122 131
rect 141 127 165 131
rect 105 126 145 127
rect 105 124 119 126
rect 121 124 145 126
rect 105 123 145 124
rect 105 112 109 123
rect 153 122 157 124
rect 161 123 167 127
rect 153 120 154 122
rect 156 120 157 122
rect 153 119 157 120
rect 153 115 160 119
rect 103 110 109 112
rect 103 108 104 110
rect 106 108 109 110
rect 103 106 109 108
rect 113 110 117 115
rect 113 108 114 110
rect 116 108 117 110
rect 113 106 117 108
rect 105 103 109 106
rect 105 99 125 103
rect 121 95 125 99
rect 156 104 160 115
rect 163 113 167 123
rect 163 111 164 113
rect 166 111 167 113
rect 163 109 167 111
rect 156 103 174 104
rect 136 101 140 103
rect 156 102 170 103
rect 136 99 137 101
rect 139 99 140 101
rect 121 94 131 95
rect 121 92 127 94
rect 129 92 131 94
rect 121 91 131 92
rect 136 94 140 99
rect 145 101 170 102
rect 172 101 174 103
rect 145 99 147 101
rect 149 100 174 101
rect 149 99 160 100
rect 145 98 160 99
rect 199 127 203 131
rect 199 123 214 127
rect 189 114 195 115
rect 210 110 214 123
rect 217 120 218 131
rect 210 108 211 110
rect 213 108 214 110
rect 210 102 214 108
rect 196 101 214 102
rect 196 99 198 101
rect 200 99 214 101
rect 196 98 214 99
rect 136 92 137 94
rect 139 93 161 94
rect 139 92 157 93
rect 136 91 157 92
rect 159 91 161 93
rect 27 90 52 91
rect 136 90 161 91
rect 166 90 170 92
rect 18 88 19 90
rect 21 88 22 90
rect 166 88 167 90
rect 169 88 170 90
rect 18 85 22 88
rect 74 87 80 88
rect 74 85 76 87
rect 78 85 80 87
rect 108 87 114 88
rect 108 85 110 87
rect 112 85 114 87
rect 166 85 170 88
rect 186 88 192 89
rect 186 86 188 88
rect 190 86 192 88
rect 186 85 192 86
rect 205 88 211 89
rect 205 86 207 88
rect 209 86 211 88
rect 205 85 211 86
rect 18 66 22 69
rect 74 67 76 69
rect 78 67 80 69
rect 74 66 80 67
rect 108 67 110 69
rect 112 67 114 69
rect 108 66 114 67
rect 166 66 170 69
rect 18 64 19 66
rect 21 64 22 66
rect 166 64 167 66
rect 169 64 170 66
rect 186 68 192 69
rect 186 66 188 68
rect 190 66 192 68
rect 186 65 192 66
rect 205 68 211 69
rect 205 66 207 68
rect 209 66 211 68
rect 205 65 211 66
rect 18 62 22 64
rect 27 63 52 64
rect 136 63 161 64
rect 27 61 29 63
rect 31 62 52 63
rect 31 61 49 62
rect 27 60 49 61
rect 51 60 52 62
rect 28 55 43 56
rect 28 54 39 55
rect 14 53 39 54
rect 41 53 43 55
rect 14 51 16 53
rect 18 52 43 53
rect 48 55 52 60
rect 57 62 67 63
rect 57 60 59 62
rect 61 60 67 62
rect 57 59 67 60
rect 48 53 49 55
rect 51 53 52 55
rect 18 51 32 52
rect 48 51 52 53
rect 14 50 32 51
rect 21 43 25 45
rect 21 41 22 43
rect 24 41 25 43
rect 21 31 25 41
rect 28 39 32 50
rect 63 55 67 59
rect 63 51 83 55
rect 79 48 83 51
rect 71 46 75 48
rect 71 44 72 46
rect 74 44 75 46
rect 71 39 75 44
rect 79 46 85 48
rect 79 44 82 46
rect 84 44 85 46
rect 79 42 85 44
rect 28 35 35 39
rect 31 34 35 35
rect 31 32 32 34
rect 34 32 35 34
rect 21 27 27 31
rect 31 30 35 32
rect 79 31 83 42
rect 43 30 83 31
rect 43 28 67 30
rect 69 28 83 30
rect 43 27 83 28
rect 23 23 47 27
rect 66 23 70 27
rect 121 62 131 63
rect 121 60 127 62
rect 129 60 131 62
rect 121 59 131 60
rect 136 62 157 63
rect 136 60 137 62
rect 139 61 157 62
rect 159 61 161 63
rect 166 62 170 64
rect 139 60 161 61
rect 121 55 125 59
rect 105 51 125 55
rect 105 48 109 51
rect 103 46 109 48
rect 103 44 104 46
rect 106 44 109 46
rect 103 42 109 44
rect 105 31 109 42
rect 113 46 117 48
rect 136 55 140 60
rect 136 53 137 55
rect 139 53 140 55
rect 136 51 140 53
rect 145 55 160 56
rect 145 53 147 55
rect 149 54 160 55
rect 149 53 174 54
rect 145 52 170 53
rect 156 51 170 52
rect 172 51 174 53
rect 156 50 174 51
rect 113 44 114 46
rect 116 44 117 46
rect 113 39 117 44
rect 156 39 160 50
rect 153 35 160 39
rect 163 43 167 45
rect 163 41 164 43
rect 166 41 167 43
rect 153 34 157 35
rect 153 32 154 34
rect 156 32 157 34
rect 105 30 145 31
rect 153 30 157 32
rect 163 31 167 41
rect 196 55 214 56
rect 196 53 198 55
rect 200 53 214 55
rect 196 52 214 53
rect 210 46 214 52
rect 210 44 211 46
rect 213 44 214 46
rect 189 39 195 40
rect 105 28 119 30
rect 121 28 145 30
rect 105 27 145 28
rect 161 27 167 31
rect 118 23 122 27
rect 141 23 165 27
rect 210 31 214 44
rect 199 27 214 31
rect 199 23 203 27
rect 217 23 218 34
rect 53 22 59 23
rect 53 20 55 22
rect 57 20 59 22
rect 18 15 24 16
rect 18 13 20 15
rect 22 13 24 15
rect 53 15 59 20
rect 66 21 67 23
rect 69 21 70 23
rect 66 19 70 21
rect 75 22 81 23
rect 75 20 77 22
rect 79 20 81 22
rect 53 13 55 15
rect 57 13 59 15
rect 75 15 81 20
rect 75 13 77 15
rect 79 13 81 15
rect 107 22 113 23
rect 107 20 109 22
rect 111 20 113 22
rect 107 15 113 20
rect 118 21 119 23
rect 121 21 122 23
rect 118 19 122 21
rect 129 22 135 23
rect 129 20 131 22
rect 133 20 135 22
rect 107 13 109 15
rect 111 13 113 15
rect 129 15 135 20
rect 186 22 203 23
rect 186 20 188 22
rect 190 20 203 22
rect 186 19 203 20
rect 129 13 131 15
rect 133 13 135 15
rect 164 15 170 16
rect 164 13 166 15
rect 168 13 170 15
rect 205 15 211 16
rect 205 13 207 15
rect 209 13 211 15
rect 18 -5 20 -3
rect 22 -5 24 -3
rect 18 -6 24 -5
rect 53 -5 55 -3
rect 57 -5 59 -3
rect 53 -10 59 -5
rect 75 -5 77 -3
rect 79 -5 81 -3
rect 53 -12 55 -10
rect 57 -12 59 -10
rect 53 -13 59 -12
rect 66 -11 70 -9
rect 66 -13 67 -11
rect 69 -13 70 -11
rect 75 -10 81 -5
rect 75 -12 77 -10
rect 79 -12 81 -10
rect 75 -13 81 -12
rect 107 -5 109 -3
rect 111 -5 113 -3
rect 107 -10 113 -5
rect 129 -5 131 -3
rect 133 -5 135 -3
rect 107 -12 109 -10
rect 111 -12 113 -10
rect 107 -13 113 -12
rect 118 -11 122 -9
rect 118 -13 119 -11
rect 121 -13 122 -11
rect 129 -10 135 -5
rect 164 -5 166 -3
rect 168 -5 170 -3
rect 164 -6 170 -5
rect 205 -5 207 -3
rect 209 -5 211 -3
rect 205 -6 211 -5
rect 129 -12 131 -10
rect 133 -12 135 -10
rect 129 -13 135 -12
rect 186 -10 203 -9
rect 186 -12 188 -10
rect 190 -12 203 -10
rect 186 -13 203 -12
rect 23 -17 47 -13
rect 66 -17 70 -13
rect 21 -21 27 -17
rect 43 -18 83 -17
rect 43 -20 67 -18
rect 69 -20 83 -18
rect 21 -31 25 -21
rect 31 -22 35 -20
rect 43 -21 83 -20
rect 31 -24 32 -22
rect 34 -24 35 -22
rect 31 -25 35 -24
rect 21 -33 22 -31
rect 24 -33 25 -31
rect 21 -35 25 -33
rect 28 -29 35 -25
rect 28 -40 32 -29
rect 71 -34 75 -29
rect 71 -36 72 -34
rect 74 -36 75 -34
rect 14 -41 32 -40
rect 14 -43 16 -41
rect 18 -42 32 -41
rect 18 -43 43 -42
rect 14 -44 39 -43
rect 28 -45 39 -44
rect 41 -45 43 -43
rect 28 -46 43 -45
rect 48 -43 52 -41
rect 48 -45 49 -43
rect 51 -45 52 -43
rect 48 -50 52 -45
rect 71 -38 75 -36
rect 79 -32 83 -21
rect 79 -34 85 -32
rect 79 -36 82 -34
rect 84 -36 85 -34
rect 79 -38 85 -36
rect 79 -41 83 -38
rect 63 -45 83 -41
rect 63 -49 67 -45
rect 27 -51 49 -50
rect 18 -54 22 -52
rect 27 -53 29 -51
rect 31 -52 49 -51
rect 51 -52 52 -50
rect 31 -53 52 -52
rect 57 -50 67 -49
rect 57 -52 59 -50
rect 61 -52 67 -50
rect 57 -53 67 -52
rect 118 -17 122 -13
rect 141 -17 165 -13
rect 105 -18 145 -17
rect 105 -20 119 -18
rect 121 -20 145 -18
rect 105 -21 145 -20
rect 105 -32 109 -21
rect 153 -22 157 -20
rect 161 -21 167 -17
rect 153 -24 154 -22
rect 156 -24 157 -22
rect 153 -25 157 -24
rect 153 -29 160 -25
rect 103 -34 109 -32
rect 103 -36 104 -34
rect 106 -36 109 -34
rect 103 -38 109 -36
rect 113 -34 117 -29
rect 113 -36 114 -34
rect 116 -36 117 -34
rect 113 -38 117 -36
rect 105 -41 109 -38
rect 105 -45 125 -41
rect 121 -49 125 -45
rect 156 -40 160 -29
rect 163 -31 167 -21
rect 163 -33 164 -31
rect 166 -33 167 -31
rect 163 -35 167 -33
rect 156 -41 174 -40
rect 136 -43 140 -41
rect 156 -42 170 -41
rect 136 -45 137 -43
rect 139 -45 140 -43
rect 121 -50 131 -49
rect 121 -52 127 -50
rect 129 -52 131 -50
rect 121 -53 131 -52
rect 136 -50 140 -45
rect 145 -43 170 -42
rect 172 -43 174 -41
rect 145 -45 147 -43
rect 149 -44 174 -43
rect 149 -45 160 -44
rect 145 -46 160 -45
rect 199 -17 203 -13
rect 199 -21 214 -17
rect 189 -30 195 -29
rect 210 -34 214 -21
rect 217 -24 218 -13
rect 210 -36 211 -34
rect 213 -36 214 -34
rect 210 -42 214 -36
rect 196 -43 214 -42
rect 196 -45 198 -43
rect 200 -45 214 -43
rect 196 -46 214 -45
rect 136 -52 137 -50
rect 139 -51 161 -50
rect 139 -52 157 -51
rect 136 -53 157 -52
rect 159 -53 161 -51
rect 27 -54 52 -53
rect 136 -54 161 -53
rect 166 -54 170 -52
rect 18 -56 19 -54
rect 21 -56 22 -54
rect 166 -56 167 -54
rect 169 -56 170 -54
rect 18 -59 22 -56
rect 74 -57 80 -56
rect 74 -59 76 -57
rect 78 -59 80 -57
rect 108 -57 114 -56
rect 108 -59 110 -57
rect 112 -59 114 -57
rect 166 -59 170 -56
rect 186 -56 192 -55
rect 186 -58 188 -56
rect 190 -58 192 -56
rect 186 -59 192 -58
rect 205 -56 211 -55
rect 205 -58 207 -56
rect 209 -58 211 -56
rect 205 -59 211 -58
rect 18 -78 22 -75
rect 74 -77 76 -75
rect 78 -77 80 -75
rect 74 -78 80 -77
rect 108 -77 110 -75
rect 112 -77 114 -75
rect 108 -78 114 -77
rect 166 -78 170 -75
rect 18 -80 19 -78
rect 21 -80 22 -78
rect 166 -80 167 -78
rect 169 -80 170 -78
rect 186 -76 192 -75
rect 186 -78 188 -76
rect 190 -78 192 -76
rect 186 -79 192 -78
rect 205 -76 211 -75
rect 205 -78 207 -76
rect 209 -78 211 -76
rect 205 -79 211 -78
rect 18 -82 22 -80
rect 27 -81 52 -80
rect 136 -81 161 -80
rect 27 -83 29 -81
rect 31 -82 52 -81
rect 31 -83 49 -82
rect 27 -84 49 -83
rect 51 -84 52 -82
rect 28 -89 43 -88
rect 28 -90 39 -89
rect 14 -91 39 -90
rect 41 -91 43 -89
rect 14 -93 16 -91
rect 18 -92 43 -91
rect 48 -89 52 -84
rect 57 -82 67 -81
rect 57 -84 59 -82
rect 61 -84 67 -82
rect 57 -85 67 -84
rect 48 -91 49 -89
rect 51 -91 52 -89
rect 18 -93 32 -92
rect 48 -93 52 -91
rect 14 -94 32 -93
rect 21 -101 25 -99
rect 21 -103 22 -101
rect 24 -103 25 -101
rect 21 -113 25 -103
rect 28 -105 32 -94
rect 63 -89 67 -85
rect 63 -93 83 -89
rect 79 -96 83 -93
rect 71 -98 75 -96
rect 71 -100 72 -98
rect 74 -100 75 -98
rect 71 -105 75 -100
rect 79 -98 85 -96
rect 79 -100 82 -98
rect 84 -100 85 -98
rect 79 -102 85 -100
rect 28 -109 35 -105
rect 31 -110 35 -109
rect 31 -112 32 -110
rect 34 -112 35 -110
rect 21 -117 27 -113
rect 31 -114 35 -112
rect 79 -113 83 -102
rect 43 -114 83 -113
rect 43 -116 67 -114
rect 69 -116 83 -114
rect 43 -117 83 -116
rect 23 -121 47 -117
rect 66 -121 70 -117
rect 121 -82 131 -81
rect 121 -84 127 -82
rect 129 -84 131 -82
rect 121 -85 131 -84
rect 136 -82 157 -81
rect 136 -84 137 -82
rect 139 -83 157 -82
rect 159 -83 161 -81
rect 166 -82 170 -80
rect 139 -84 161 -83
rect 121 -89 125 -85
rect 105 -93 125 -89
rect 105 -96 109 -93
rect 103 -98 109 -96
rect 103 -100 104 -98
rect 106 -100 109 -98
rect 103 -102 109 -100
rect 105 -113 109 -102
rect 113 -98 117 -96
rect 136 -89 140 -84
rect 136 -91 137 -89
rect 139 -91 140 -89
rect 136 -93 140 -91
rect 145 -89 160 -88
rect 145 -91 147 -89
rect 149 -90 160 -89
rect 149 -91 174 -90
rect 145 -92 170 -91
rect 156 -93 170 -92
rect 172 -93 174 -91
rect 156 -94 174 -93
rect 113 -100 114 -98
rect 116 -100 117 -98
rect 113 -105 117 -100
rect 156 -105 160 -94
rect 153 -109 160 -105
rect 163 -101 167 -99
rect 163 -103 164 -101
rect 166 -103 167 -101
rect 153 -110 157 -109
rect 153 -112 154 -110
rect 156 -112 157 -110
rect 105 -114 145 -113
rect 153 -114 157 -112
rect 163 -113 167 -103
rect 196 -89 214 -88
rect 196 -91 198 -89
rect 200 -91 214 -89
rect 196 -92 214 -91
rect 210 -98 214 -92
rect 210 -100 211 -98
rect 213 -100 214 -98
rect 189 -105 195 -104
rect 105 -116 119 -114
rect 121 -116 145 -114
rect 105 -117 145 -116
rect 161 -117 167 -113
rect 118 -121 122 -117
rect 141 -121 165 -117
rect 210 -113 214 -100
rect 199 -117 214 -113
rect 199 -121 203 -117
rect 217 -121 218 -110
rect 53 -122 59 -121
rect 53 -124 55 -122
rect 57 -124 59 -122
rect 18 -129 24 -128
rect 18 -131 20 -129
rect 22 -131 24 -129
rect 53 -129 59 -124
rect 66 -123 67 -121
rect 69 -123 70 -121
rect 66 -125 70 -123
rect 75 -122 81 -121
rect 75 -124 77 -122
rect 79 -124 81 -122
rect 53 -131 55 -129
rect 57 -131 59 -129
rect 75 -129 81 -124
rect 75 -131 77 -129
rect 79 -131 81 -129
rect 107 -122 113 -121
rect 107 -124 109 -122
rect 111 -124 113 -122
rect 107 -129 113 -124
rect 118 -123 119 -121
rect 121 -123 122 -121
rect 118 -125 122 -123
rect 129 -122 135 -121
rect 129 -124 131 -122
rect 133 -124 135 -122
rect 107 -131 109 -129
rect 111 -131 113 -129
rect 129 -129 135 -124
rect 186 -122 203 -121
rect 186 -124 188 -122
rect 190 -124 203 -122
rect 186 -125 203 -124
rect 129 -131 131 -129
rect 133 -131 135 -129
rect 164 -129 170 -128
rect 164 -131 166 -129
rect 168 -131 170 -129
rect 205 -129 211 -128
rect 205 -131 207 -129
rect 209 -131 211 -129
<< via1 >>
rect 8 100 10 102
rect 89 108 91 110
rect 99 121 101 123
rect 130 100 132 102
rect 187 121 189 123
rect 187 108 189 110
rect 219 104 221 106
rect 8 52 10 54
rect 89 44 91 46
rect 130 52 132 54
rect 99 31 101 33
rect 147 39 149 41
rect 187 50 189 52
rect 187 31 189 33
rect 211 20 213 22
rect 8 -44 10 -42
rect 89 -36 91 -34
rect 99 -23 101 -21
rect 147 -28 149 -26
rect 130 -44 132 -42
rect 187 -19 189 -17
rect 187 -36 189 -34
rect 219 -40 221 -38
rect 8 -92 10 -90
rect 89 -100 91 -98
rect 130 -92 132 -90
rect 99 -113 101 -111
rect 147 -105 149 -103
rect 187 -94 189 -92
rect 187 -113 189 -111
<< via2 >>
rect 223 104 225 106
rect 223 39 225 41
rect 223 -40 225 -38
rect 223 -105 225 -103
<< labels >>
rlabel alu1 53 81 53 81 1 gnd
rlabel alu1 135 81 135 81 1 gnd
rlabel alu1 132 117 132 117 1 cin
rlabel alu1 135 73 135 73 5 gnd
rlabel alu1 53 73 53 73 5 gnd
rlabel alu1 57 117 57 117 1 b_0
rlabel alu1 65 109 65 109 1 a_0
rlabel alu1 65 45 65 45 1 a_1
rlabel alu1 57 37 57 37 1 b_1
rlabel alu1 179 45 179 45 1 s_1
rlabel alu1 179 114 179 114 1 s_0
rlabel alu1 158 145 158 145 1 Vdd
rlabel alu1 184 145 184 145 1 Vdd
rlabel alu1 94 145 94 145 1 Vdd
rlabel alu1 29 145 29 145 1 vdd
rlabel alu1 29 8 29 8 1 Vdd
rlabel alu1 94 9 94 9 1 Vdd
rlabel alu1 185 9 185 9 1 Vdd
rlabel alu1 159 9 159 9 1 Vdd
rlabel alu1 159 -135 159 -135 1 Vdd
rlabel alu1 185 -135 185 -135 1 Vdd
rlabel alu1 94 -135 94 -135 1 Vdd
rlabel alu1 29 -136 29 -136 1 Vdd
rlabel alu1 29 1 29 1 1 vdd
rlabel alu1 94 1 94 1 1 Vdd
rlabel alu1 184 1 184 1 1 Vdd
rlabel alu1 158 1 158 1 1 Vdd
rlabel alu1 53 -71 53 -71 5 gnd
rlabel alu1 135 -71 135 -71 5 gnd
rlabel alu1 220 -105 220 -105 5 cout
rlabel alu1 135 -63 135 -63 1 gnd
rlabel alu1 53 -63 53 -63 1 gnd
rlabel alu1 179 -30 179 -30 1 s_2
rlabel alu1 179 -99 179 -99 1 s_3
rlabel alu1 57 -107 57 -107 1 b_3
rlabel alu1 65 -99 65 -99 1 a_3
rlabel alu1 57 -27 57 -27 1 b_2
rlabel alu1 65 -35 65 -35 1 a_2
<< end >>
