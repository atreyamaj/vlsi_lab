magic
tech scmos
timestamp 1520960406
<< nwell >>
rect -24 10 36 27
<< polysilicon >>
rect -21 21 -19 24
rect -8 21 -6 24
rect 18 21 20 24
rect -21 2 -19 15
rect -8 2 -6 15
rect 18 2 20 15
rect -20 -2 -19 2
rect -7 -2 -6 2
rect 19 -2 20 2
rect -21 -9 -19 -2
rect -8 -9 -6 -2
rect 18 -12 20 -2
rect -21 -18 -19 -15
rect -8 -18 -6 -15
rect 18 -18 20 -15
<< ndiffusion >>
rect -24 -10 -21 -9
rect -22 -14 -21 -10
rect -24 -15 -21 -14
rect -19 -15 -8 -9
rect -6 -10 -2 -9
rect -6 -14 -4 -10
rect -6 -15 -2 -14
rect 9 -15 18 -12
rect 20 -15 30 -12
<< pdiffusion >>
rect -24 20 -21 21
rect -22 16 -21 20
rect -24 15 -21 16
rect -19 20 -8 21
rect -19 16 -16 20
rect -12 16 -8 20
rect -19 15 -8 16
rect -6 20 -2 21
rect 6 20 18 21
rect -6 16 -4 20
rect 9 16 18 20
rect -6 15 -2 16
rect 6 15 18 16
rect 20 20 33 21
rect 20 16 30 20
rect 20 15 33 16
<< metal1 >>
rect -26 29 36 30
rect -26 27 -3 29
rect -16 20 -13 27
rect 1 27 36 29
rect 6 20 9 27
rect 34 16 35 19
rect -26 8 -23 16
rect -3 8 0 16
rect -26 5 0 8
rect -3 1 0 5
rect -3 -2 15 1
rect -3 -10 0 -2
rect 32 -11 35 16
rect -26 -21 -23 -14
rect 34 -14 35 -11
rect 5 -21 8 -15
rect -26 -24 36 -21
<< ntransistor >>
rect -21 -15 -19 -9
rect -8 -15 -6 -9
rect 18 -15 20 -12
<< ptransistor >>
rect -21 15 -19 21
rect -8 15 -6 21
rect 18 15 20 21
<< polycontact >>
rect -24 -2 -20 2
rect -11 -2 -7 2
rect 15 -2 19 2
<< ndcontact >>
rect -26 -14 -22 -10
rect -4 -14 0 -10
rect 5 -15 9 -11
rect 30 -15 34 -11
<< pdcontact >>
rect -26 16 -22 20
rect -16 16 -12 20
rect -4 16 0 20
rect 5 16 9 20
rect 30 16 34 20
<< nsubstratencontact >>
rect -3 25 1 29
<< labels >>
rlabel polycontact -22 0 -22 0 3 A
rlabel polycontact -9 0 -9 0 1 B
rlabel metal1 8 29 8 29 5 vdd
rlabel ndiffusion -16 -12 -16 -12 1 n1
rlabel metal1 7 0 7 0 1 nand_out
rlabel metal1 34 -2 34 -2 7 out
rlabel metal1 6 -23 6 -23 1 gnd
<< end >>
