* SPICE3 file created from nand.ext - technology: scmos

.include /home/vlsilab/UG_students_2018/t14y_tsmc_025_level3.txt

M1000 out A vdd vdd cmosp w=8u l=2u
+  ad=56p pd=30u as=80p ps=52u
M1001 vdd B out vdd cmosp w=8u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1002 n1 A out Gnd cmosn w=4u l=2u
+  ad=28p pd=22u as=20p ps=18u
M1003 gnd B n1 Gnd cmosn w=4u l=2u
+  ad=28p pd=22u as=0p ps=0u
C0 out Gnd 2.54fF
C1 B Gnd 4.76fF
C2 A Gnd 7.30fF
C3 vdd Gnd 3.10fF

gd gnd 0 0
v_dd vdd 0 3.3

vin_a A 0 PULSE(0 3.3 0ns 0.1ns 0.1ns 2us 4.2us)
vin_b B 0 PULSE(0 3.3 0ns 0.1ns 0.1ns 3us 6.2us)

.control
tran 0.1ns 20us
run
plot (out) (0.5*A) (0.25*B)
.endc

.end
