magic
tech scmos
timestamp 1553857537
<< rotate >>
rect 75 156 86 158
rect 52 152 54 154
rect 75 149 89 156
rect 78 147 89 149
rect 75 12 86 14
rect 52 8 54 10
rect 75 5 89 12
rect 78 3 89 5
<< ab >>
rect -75 279 182 293
rect -75 275 7 279
rect 9 275 179 279
rect 181 275 182 279
rect -75 167 182 275
rect -75 163 7 167
rect 9 163 179 167
rect 181 163 182 167
rect -75 135 182 163
rect -75 131 7 135
rect 9 131 179 135
rect 181 131 182 135
rect -75 23 182 131
rect -75 19 7 23
rect 9 19 179 23
rect 181 19 182 23
rect -75 5 182 19
rect 184 182 225 293
rect 184 179 226 182
rect 184 38 225 179
rect 184 35 226 38
rect 184 5 225 35
<< nwell >>
rect -80 253 228 298
rect -80 109 228 189
rect -80 0 228 45
<< pwell >>
rect -80 189 228 253
rect -80 45 228 109
<< poly >>
rect -66 280 -64 285
rect -56 280 -54 285
rect 14 287 16 291
rect -46 278 -44 282
rect -26 280 -24 285
rect -16 280 -14 285
rect -66 264 -64 267
rect -70 262 -64 264
rect -70 260 -68 262
rect -66 260 -64 262
rect -70 258 -64 260
rect -66 245 -64 258
rect -56 256 -54 267
rect -6 278 -4 282
rect -26 264 -24 267
rect -30 262 -24 264
rect -30 260 -28 262
rect -26 260 -24 262
rect -46 256 -44 260
rect -30 258 -24 260
rect -60 254 -54 256
rect -60 252 -58 254
rect -56 252 -54 254
rect -60 250 -54 252
rect -50 254 -44 256
rect -50 252 -48 254
rect -46 252 -44 254
rect -50 250 -44 252
rect -59 245 -57 250
rect -46 245 -44 250
rect -26 245 -24 258
rect -16 256 -14 267
rect 37 284 39 289
rect 44 284 46 289
rect 62 287 64 291
rect 72 287 74 291
rect 82 287 84 291
rect 104 287 106 291
rect 114 287 116 291
rect 124 287 126 291
rect 27 275 29 280
rect -6 256 -4 260
rect -20 254 -14 256
rect -20 252 -18 254
rect -16 252 -14 254
rect -20 250 -14 252
rect -10 254 -4 256
rect -10 252 -8 254
rect -6 252 -4 254
rect -10 250 -4 252
rect -19 245 -17 250
rect -6 245 -4 250
rect 14 249 16 262
rect 27 259 29 262
rect 142 284 144 289
rect 149 284 151 289
rect 172 287 174 291
rect 193 287 195 291
rect 200 287 202 291
rect 159 275 161 280
rect 213 277 215 282
rect 193 263 195 266
rect 159 259 161 262
rect 20 257 29 259
rect 20 255 22 257
rect 24 255 26 257
rect 37 256 39 259
rect 44 256 46 259
rect 62 256 64 259
rect 72 256 74 259
rect 82 256 84 259
rect 104 256 106 259
rect 114 256 116 259
rect 124 256 126 259
rect 142 256 144 259
rect 149 256 151 259
rect 159 257 168 259
rect 20 253 26 255
rect 14 247 20 249
rect 14 245 16 247
rect 18 245 20 247
rect -66 229 -64 234
rect -59 229 -57 234
rect -46 232 -44 236
rect 14 243 20 245
rect 14 240 16 243
rect 24 240 26 253
rect 34 254 40 256
rect 34 252 36 254
rect 38 252 40 254
rect 34 250 40 252
rect 44 254 66 256
rect 44 252 55 254
rect 57 252 62 254
rect 64 252 66 254
rect 44 250 66 252
rect 70 254 76 256
rect 70 252 72 254
rect 74 252 76 254
rect 70 250 76 252
rect 80 254 86 256
rect 80 252 82 254
rect 84 252 86 254
rect 80 250 86 252
rect 102 254 108 256
rect 102 252 104 254
rect 106 252 108 254
rect 102 250 108 252
rect 112 254 118 256
rect 112 252 114 254
rect 116 252 118 254
rect 112 250 118 252
rect 122 254 144 256
rect 122 252 124 254
rect 126 252 131 254
rect 133 252 144 254
rect 122 250 144 252
rect 148 254 154 256
rect 148 252 150 254
rect 152 252 154 254
rect 148 250 154 252
rect 34 247 36 250
rect 44 247 46 250
rect 64 247 66 250
rect 71 247 73 250
rect -26 229 -24 234
rect -19 229 -17 234
rect -6 232 -4 236
rect 14 223 16 227
rect 24 225 26 230
rect 34 228 36 233
rect 44 228 46 233
rect 82 241 84 250
rect 104 241 106 250
rect 115 247 117 250
rect 122 247 124 250
rect 142 247 144 250
rect 152 247 154 250
rect 162 255 164 257
rect 166 255 168 257
rect 162 253 168 255
rect 162 240 164 253
rect 172 249 174 262
rect 189 261 195 263
rect 189 259 191 261
rect 193 259 195 261
rect 189 257 195 259
rect 168 247 174 249
rect 193 247 195 257
rect 200 256 202 266
rect 213 256 215 259
rect 199 254 205 256
rect 199 252 201 254
rect 203 252 205 254
rect 199 250 205 252
rect 209 254 215 256
rect 209 252 211 254
rect 213 252 215 254
rect 209 250 215 252
rect 203 247 205 250
rect 213 247 215 250
rect 168 245 170 247
rect 172 245 174 247
rect 168 243 174 245
rect 172 240 174 243
rect 142 228 144 233
rect 152 228 154 233
rect 64 223 66 227
rect 71 223 73 227
rect 82 223 84 227
rect 104 223 106 227
rect 115 223 117 227
rect 122 223 124 227
rect 162 225 164 230
rect 193 236 195 241
rect 203 236 205 241
rect 213 233 215 238
rect 172 223 174 227
rect -66 208 -64 213
rect -59 208 -57 213
rect -46 206 -44 210
rect -26 208 -24 213
rect -19 208 -17 213
rect 14 215 16 219
rect -6 206 -4 210
rect 24 212 26 217
rect 64 215 66 219
rect 71 215 73 219
rect 82 215 84 219
rect 104 215 106 219
rect 115 215 117 219
rect 122 215 124 219
rect 34 209 36 214
rect 44 209 46 214
rect 14 199 16 202
rect 14 197 20 199
rect -66 184 -64 197
rect -59 192 -57 197
rect -46 192 -44 197
rect -60 190 -54 192
rect -60 188 -58 190
rect -56 188 -54 190
rect -60 186 -54 188
rect -50 190 -44 192
rect -50 188 -48 190
rect -46 188 -44 190
rect -50 186 -44 188
rect -70 182 -64 184
rect -70 180 -68 182
rect -66 180 -64 182
rect -70 178 -64 180
rect -66 175 -64 178
rect -56 175 -54 186
rect -46 182 -44 186
rect -26 184 -24 197
rect -19 192 -17 197
rect -6 192 -4 197
rect -20 190 -14 192
rect -20 188 -18 190
rect -16 188 -14 190
rect -20 186 -14 188
rect -10 190 -4 192
rect -10 188 -8 190
rect -6 188 -4 190
rect -10 186 -4 188
rect -30 182 -24 184
rect -30 180 -28 182
rect -26 180 -24 182
rect -30 178 -24 180
rect -26 175 -24 178
rect -16 175 -14 186
rect -6 182 -4 186
rect 14 195 16 197
rect 18 195 20 197
rect 14 193 20 195
rect -66 157 -64 162
rect -56 157 -54 162
rect -46 160 -44 164
rect 14 180 16 193
rect 24 189 26 202
rect 20 187 26 189
rect 20 185 22 187
rect 24 185 26 187
rect 34 192 36 195
rect 44 192 46 195
rect 64 192 66 195
rect 71 192 73 195
rect 82 192 84 201
rect 104 192 106 201
rect 142 209 144 214
rect 152 209 154 214
rect 162 212 164 217
rect 172 215 174 219
rect 115 192 117 195
rect 122 192 124 195
rect 142 192 144 195
rect 152 192 154 195
rect 34 190 40 192
rect 34 188 36 190
rect 38 188 40 190
rect 34 186 40 188
rect 44 190 66 192
rect 44 188 55 190
rect 57 188 62 190
rect 64 188 66 190
rect 44 186 66 188
rect 70 190 76 192
rect 70 188 72 190
rect 74 188 76 190
rect 70 186 76 188
rect 80 190 86 192
rect 80 188 82 190
rect 84 188 86 190
rect 80 186 86 188
rect 102 190 108 192
rect 102 188 104 190
rect 106 188 108 190
rect 102 186 108 188
rect 112 190 118 192
rect 112 188 114 190
rect 116 188 118 190
rect 112 186 118 188
rect 122 190 144 192
rect 122 188 124 190
rect 126 188 131 190
rect 133 188 144 190
rect 122 186 144 188
rect 148 190 154 192
rect 148 188 150 190
rect 152 188 154 190
rect 148 186 154 188
rect 162 189 164 202
rect 172 199 174 202
rect 168 197 174 199
rect 168 195 170 197
rect 172 195 174 197
rect 193 201 195 206
rect 203 201 205 206
rect 213 204 215 209
rect 168 193 174 195
rect 162 187 168 189
rect 20 183 29 185
rect 37 183 39 186
rect 44 183 46 186
rect 62 183 64 186
rect 72 183 74 186
rect 82 183 84 186
rect 104 183 106 186
rect 114 183 116 186
rect 124 183 126 186
rect 142 183 144 186
rect 149 183 151 186
rect 162 185 164 187
rect 166 185 168 187
rect 159 183 168 185
rect 27 180 29 183
rect -26 157 -24 162
rect -16 157 -14 162
rect -6 160 -4 164
rect 27 162 29 167
rect 14 151 16 155
rect 37 153 39 158
rect 44 153 46 158
rect 159 180 161 183
rect 172 180 174 193
rect 193 185 195 195
rect 203 192 205 195
rect 213 192 215 195
rect 199 190 205 192
rect 199 188 201 190
rect 203 188 205 190
rect 199 186 205 188
rect 209 190 215 192
rect 209 188 211 190
rect 213 188 215 190
rect 209 186 215 188
rect 189 183 195 185
rect 189 181 191 183
rect 193 181 195 183
rect 159 162 161 167
rect 62 151 64 155
rect 72 151 74 155
rect 82 151 84 155
rect 104 151 106 155
rect 114 151 116 155
rect 124 151 126 155
rect 142 153 144 158
rect 149 153 151 158
rect 189 179 195 181
rect 193 176 195 179
rect 200 176 202 186
rect 213 183 215 186
rect 213 160 215 165
rect 172 151 174 155
rect 193 151 195 155
rect 200 151 202 155
rect -66 136 -64 141
rect -56 136 -54 141
rect 14 143 16 147
rect -46 134 -44 138
rect -26 136 -24 141
rect -16 136 -14 141
rect -66 120 -64 123
rect -70 118 -64 120
rect -70 116 -68 118
rect -66 116 -64 118
rect -70 114 -64 116
rect -66 101 -64 114
rect -56 112 -54 123
rect -6 134 -4 138
rect -26 120 -24 123
rect -30 118 -24 120
rect -30 116 -28 118
rect -26 116 -24 118
rect -46 112 -44 116
rect -30 114 -24 116
rect -60 110 -54 112
rect -60 108 -58 110
rect -56 108 -54 110
rect -60 106 -54 108
rect -50 110 -44 112
rect -50 108 -48 110
rect -46 108 -44 110
rect -50 106 -44 108
rect -59 101 -57 106
rect -46 101 -44 106
rect -26 101 -24 114
rect -16 112 -14 123
rect 37 140 39 145
rect 44 140 46 145
rect 62 143 64 147
rect 72 143 74 147
rect 82 143 84 147
rect 104 143 106 147
rect 114 143 116 147
rect 124 143 126 147
rect 27 131 29 136
rect -6 112 -4 116
rect -20 110 -14 112
rect -20 108 -18 110
rect -16 108 -14 110
rect -20 106 -14 108
rect -10 110 -4 112
rect -10 108 -8 110
rect -6 108 -4 110
rect -10 106 -4 108
rect -19 101 -17 106
rect -6 101 -4 106
rect 14 105 16 118
rect 27 115 29 118
rect 142 140 144 145
rect 149 140 151 145
rect 172 143 174 147
rect 193 143 195 147
rect 200 143 202 147
rect 159 131 161 136
rect 213 133 215 138
rect 193 119 195 122
rect 159 115 161 118
rect 20 113 29 115
rect 20 111 22 113
rect 24 111 26 113
rect 37 112 39 115
rect 44 112 46 115
rect 62 112 64 115
rect 72 112 74 115
rect 82 112 84 115
rect 104 112 106 115
rect 114 112 116 115
rect 124 112 126 115
rect 142 112 144 115
rect 149 112 151 115
rect 159 113 168 115
rect 20 109 26 111
rect 14 103 20 105
rect 14 101 16 103
rect 18 101 20 103
rect -66 85 -64 90
rect -59 85 -57 90
rect -46 88 -44 92
rect 14 99 20 101
rect 14 96 16 99
rect 24 96 26 109
rect 34 110 40 112
rect 34 108 36 110
rect 38 108 40 110
rect 34 106 40 108
rect 44 110 66 112
rect 44 108 55 110
rect 57 108 62 110
rect 64 108 66 110
rect 44 106 66 108
rect 70 110 76 112
rect 70 108 72 110
rect 74 108 76 110
rect 70 106 76 108
rect 80 110 86 112
rect 80 108 82 110
rect 84 108 86 110
rect 80 106 86 108
rect 102 110 108 112
rect 102 108 104 110
rect 106 108 108 110
rect 102 106 108 108
rect 112 110 118 112
rect 112 108 114 110
rect 116 108 118 110
rect 112 106 118 108
rect 122 110 144 112
rect 122 108 124 110
rect 126 108 131 110
rect 133 108 144 110
rect 122 106 144 108
rect 148 110 154 112
rect 148 108 150 110
rect 152 108 154 110
rect 148 106 154 108
rect 34 103 36 106
rect 44 103 46 106
rect 64 103 66 106
rect 71 103 73 106
rect -26 85 -24 90
rect -19 85 -17 90
rect -6 88 -4 92
rect 14 79 16 83
rect 24 81 26 86
rect 34 84 36 89
rect 44 84 46 89
rect 82 97 84 106
rect 104 97 106 106
rect 115 103 117 106
rect 122 103 124 106
rect 142 103 144 106
rect 152 103 154 106
rect 162 111 164 113
rect 166 111 168 113
rect 162 109 168 111
rect 162 96 164 109
rect 172 105 174 118
rect 189 117 195 119
rect 189 115 191 117
rect 193 115 195 117
rect 189 113 195 115
rect 168 103 174 105
rect 193 103 195 113
rect 200 112 202 122
rect 213 112 215 115
rect 199 110 205 112
rect 199 108 201 110
rect 203 108 205 110
rect 199 106 205 108
rect 209 110 215 112
rect 209 108 211 110
rect 213 108 215 110
rect 209 106 215 108
rect 203 103 205 106
rect 213 103 215 106
rect 168 101 170 103
rect 172 101 174 103
rect 168 99 174 101
rect 172 96 174 99
rect 142 84 144 89
rect 152 84 154 89
rect 64 79 66 83
rect 71 79 73 83
rect 82 79 84 83
rect 104 79 106 83
rect 115 79 117 83
rect 122 79 124 83
rect 162 81 164 86
rect 193 92 195 97
rect 203 92 205 97
rect 213 89 215 94
rect 172 79 174 83
rect -66 64 -64 69
rect -59 64 -57 69
rect -46 62 -44 66
rect -26 64 -24 69
rect -19 64 -17 69
rect 14 71 16 75
rect -6 62 -4 66
rect 24 68 26 73
rect 64 71 66 75
rect 71 71 73 75
rect 82 71 84 75
rect 104 71 106 75
rect 115 71 117 75
rect 122 71 124 75
rect 34 65 36 70
rect 44 65 46 70
rect 14 55 16 58
rect 14 53 20 55
rect -66 40 -64 53
rect -59 48 -57 53
rect -46 48 -44 53
rect -60 46 -54 48
rect -60 44 -58 46
rect -56 44 -54 46
rect -60 42 -54 44
rect -50 46 -44 48
rect -50 44 -48 46
rect -46 44 -44 46
rect -50 42 -44 44
rect -70 38 -64 40
rect -70 36 -68 38
rect -66 36 -64 38
rect -70 34 -64 36
rect -66 31 -64 34
rect -56 31 -54 42
rect -46 38 -44 42
rect -26 40 -24 53
rect -19 48 -17 53
rect -6 48 -4 53
rect -20 46 -14 48
rect -20 44 -18 46
rect -16 44 -14 46
rect -20 42 -14 44
rect -10 46 -4 48
rect -10 44 -8 46
rect -6 44 -4 46
rect -10 42 -4 44
rect -30 38 -24 40
rect -30 36 -28 38
rect -26 36 -24 38
rect -30 34 -24 36
rect -26 31 -24 34
rect -16 31 -14 42
rect -6 38 -4 42
rect 14 51 16 53
rect 18 51 20 53
rect 14 49 20 51
rect -66 13 -64 18
rect -56 13 -54 18
rect -46 16 -44 20
rect 14 36 16 49
rect 24 45 26 58
rect 20 43 26 45
rect 20 41 22 43
rect 24 41 26 43
rect 34 48 36 51
rect 44 48 46 51
rect 64 48 66 51
rect 71 48 73 51
rect 82 48 84 57
rect 104 48 106 57
rect 142 65 144 70
rect 152 65 154 70
rect 162 68 164 73
rect 172 71 174 75
rect 115 48 117 51
rect 122 48 124 51
rect 142 48 144 51
rect 152 48 154 51
rect 34 46 40 48
rect 34 44 36 46
rect 38 44 40 46
rect 34 42 40 44
rect 44 46 66 48
rect 44 44 55 46
rect 57 44 62 46
rect 64 44 66 46
rect 44 42 66 44
rect 70 46 76 48
rect 70 44 72 46
rect 74 44 76 46
rect 70 42 76 44
rect 80 46 86 48
rect 80 44 82 46
rect 84 44 86 46
rect 80 42 86 44
rect 102 46 108 48
rect 102 44 104 46
rect 106 44 108 46
rect 102 42 108 44
rect 112 46 118 48
rect 112 44 114 46
rect 116 44 118 46
rect 112 42 118 44
rect 122 46 144 48
rect 122 44 124 46
rect 126 44 131 46
rect 133 44 144 46
rect 122 42 144 44
rect 148 46 154 48
rect 148 44 150 46
rect 152 44 154 46
rect 148 42 154 44
rect 162 45 164 58
rect 172 55 174 58
rect 168 53 174 55
rect 168 51 170 53
rect 172 51 174 53
rect 193 57 195 62
rect 203 57 205 62
rect 213 60 215 65
rect 168 49 174 51
rect 162 43 168 45
rect 20 39 29 41
rect 37 39 39 42
rect 44 39 46 42
rect 62 39 64 42
rect 72 39 74 42
rect 82 39 84 42
rect 104 39 106 42
rect 114 39 116 42
rect 124 39 126 42
rect 142 39 144 42
rect 149 39 151 42
rect 162 41 164 43
rect 166 41 168 43
rect 159 39 168 41
rect 27 36 29 39
rect -26 13 -24 18
rect -16 13 -14 18
rect -6 16 -4 20
rect 27 18 29 23
rect 14 7 16 11
rect 37 9 39 14
rect 44 9 46 14
rect 159 36 161 39
rect 172 36 174 49
rect 193 41 195 51
rect 203 48 205 51
rect 213 48 215 51
rect 199 46 205 48
rect 199 44 201 46
rect 203 44 205 46
rect 199 42 205 44
rect 209 46 215 48
rect 209 44 211 46
rect 213 44 215 46
rect 209 42 215 44
rect 189 39 195 41
rect 189 37 191 39
rect 193 37 195 39
rect 159 18 161 23
rect 62 7 64 11
rect 72 7 74 11
rect 82 7 84 11
rect 104 7 106 11
rect 114 7 116 11
rect 124 7 126 11
rect 142 9 144 14
rect 149 9 151 14
rect 189 35 195 37
rect 193 32 195 35
rect 200 32 202 42
rect 213 39 215 42
rect 213 16 215 21
rect 172 7 174 11
rect 193 7 195 11
rect 200 7 202 11
<< ndif >>
rect -71 240 -66 245
rect -73 238 -66 240
rect -73 236 -71 238
rect -69 236 -66 238
rect -73 234 -66 236
rect -64 234 -59 245
rect -57 236 -46 245
rect -44 242 -39 245
rect -44 240 -37 242
rect -31 240 -26 245
rect -44 238 -41 240
rect -39 238 -37 240
rect -44 236 -37 238
rect -33 238 -26 240
rect -33 236 -31 238
rect -29 236 -26 238
rect -57 234 -48 236
rect -55 228 -48 234
rect -33 234 -26 236
rect -24 234 -19 245
rect -17 236 -6 245
rect -4 242 1 245
rect -4 240 3 242
rect 29 240 34 247
rect -4 238 -1 240
rect 1 238 3 240
rect -4 236 3 238
rect 7 238 14 240
rect 7 236 9 238
rect 11 236 14 238
rect -17 234 -8 236
rect -55 226 -52 228
rect -50 226 -48 228
rect -55 224 -48 226
rect -15 228 -8 234
rect 7 234 14 236
rect -15 226 -12 228
rect -10 226 -8 228
rect -15 224 -8 226
rect 9 227 14 234
rect 16 234 24 240
rect 16 232 19 234
rect 21 232 24 234
rect 16 230 24 232
rect 26 237 34 240
rect 26 235 29 237
rect 31 235 34 237
rect 26 233 34 235
rect 36 245 44 247
rect 36 243 39 245
rect 41 243 44 245
rect 36 233 44 243
rect 46 245 53 247
rect 46 243 49 245
rect 51 243 53 245
rect 46 238 53 243
rect 59 240 64 247
rect 46 236 49 238
rect 51 236 53 238
rect 46 233 53 236
rect 57 238 64 240
rect 57 236 59 238
rect 61 236 64 238
rect 57 234 64 236
rect 26 230 31 233
rect 16 227 21 230
rect 59 227 64 234
rect 66 227 71 247
rect 73 241 80 247
rect 108 241 115 247
rect 73 231 82 241
rect 73 229 76 231
rect 78 229 82 231
rect 73 227 82 229
rect 84 238 91 241
rect 84 236 87 238
rect 89 236 91 238
rect 84 234 91 236
rect 97 238 104 241
rect 97 236 99 238
rect 101 236 104 238
rect 97 234 104 236
rect 84 227 89 234
rect 99 227 104 234
rect 106 231 115 241
rect 106 229 110 231
rect 112 229 115 231
rect 106 227 115 229
rect 117 227 122 247
rect 124 240 129 247
rect 135 245 142 247
rect 135 243 137 245
rect 139 243 142 245
rect 124 238 131 240
rect 124 236 127 238
rect 129 236 131 238
rect 124 234 131 236
rect 135 238 142 243
rect 135 236 137 238
rect 139 236 142 238
rect 124 227 129 234
rect 135 233 142 236
rect 144 245 152 247
rect 144 243 147 245
rect 149 243 152 245
rect 144 233 152 243
rect 154 240 159 247
rect 186 241 193 247
rect 195 245 203 247
rect 195 243 198 245
rect 200 243 203 245
rect 195 241 203 243
rect 205 241 213 247
rect 154 237 162 240
rect 154 235 157 237
rect 159 235 162 237
rect 154 233 162 235
rect 157 230 162 233
rect 164 234 172 240
rect 164 232 167 234
rect 169 232 172 234
rect 164 230 172 232
rect 167 227 172 230
rect 174 238 181 240
rect 174 236 177 238
rect 179 236 181 238
rect 174 234 181 236
rect 186 234 191 241
rect 207 238 213 241
rect 215 245 222 247
rect 215 243 218 245
rect 220 243 222 245
rect 215 241 222 243
rect 215 238 220 241
rect 207 234 211 238
rect 174 227 179 234
rect 186 232 192 234
rect 186 230 188 232
rect 190 230 192 232
rect 186 228 192 230
rect 205 232 211 234
rect 205 230 207 232
rect 209 230 211 232
rect 205 228 211 230
rect -55 216 -48 218
rect -55 214 -52 216
rect -50 214 -48 216
rect -55 208 -48 214
rect -15 216 -8 218
rect -15 214 -12 216
rect -10 214 -8 216
rect -73 206 -66 208
rect -73 204 -71 206
rect -69 204 -66 206
rect -73 202 -66 204
rect -71 197 -66 202
rect -64 197 -59 208
rect -57 206 -48 208
rect -15 208 -8 214
rect -33 206 -26 208
rect -57 197 -46 206
rect -44 204 -37 206
rect -44 202 -41 204
rect -39 202 -37 204
rect -33 204 -31 206
rect -29 204 -26 206
rect -33 202 -26 204
rect -44 200 -37 202
rect -44 197 -39 200
rect -31 197 -26 202
rect -24 197 -19 208
rect -17 206 -8 208
rect 9 208 14 215
rect 7 206 14 208
rect -17 197 -6 206
rect -4 204 3 206
rect -4 202 -1 204
rect 1 202 3 204
rect 7 204 9 206
rect 11 204 14 206
rect 7 202 14 204
rect 16 212 21 215
rect 16 210 24 212
rect 16 208 19 210
rect 21 208 24 210
rect 16 202 24 208
rect 26 209 31 212
rect 26 207 34 209
rect 26 205 29 207
rect 31 205 34 207
rect 26 202 34 205
rect -4 200 3 202
rect -4 197 1 200
rect 29 195 34 202
rect 36 199 44 209
rect 36 197 39 199
rect 41 197 44 199
rect 36 195 44 197
rect 46 206 53 209
rect 59 208 64 215
rect 46 204 49 206
rect 51 204 53 206
rect 46 199 53 204
rect 57 206 64 208
rect 57 204 59 206
rect 61 204 64 206
rect 57 202 64 204
rect 46 197 49 199
rect 51 197 53 199
rect 46 195 53 197
rect 59 195 64 202
rect 66 195 71 215
rect 73 213 82 215
rect 73 211 76 213
rect 78 211 82 213
rect 73 201 82 211
rect 84 208 89 215
rect 99 208 104 215
rect 84 206 91 208
rect 84 204 87 206
rect 89 204 91 206
rect 84 201 91 204
rect 97 206 104 208
rect 97 204 99 206
rect 101 204 104 206
rect 97 201 104 204
rect 106 213 115 215
rect 106 211 110 213
rect 112 211 115 213
rect 106 201 115 211
rect 73 195 80 201
rect 108 195 115 201
rect 117 195 122 215
rect 124 208 129 215
rect 167 212 172 215
rect 157 209 162 212
rect 124 206 131 208
rect 124 204 127 206
rect 129 204 131 206
rect 124 202 131 204
rect 135 206 142 209
rect 135 204 137 206
rect 139 204 142 206
rect 124 195 129 202
rect 135 199 142 204
rect 135 197 137 199
rect 139 197 142 199
rect 135 195 142 197
rect 144 199 152 209
rect 144 197 147 199
rect 149 197 152 199
rect 144 195 152 197
rect 154 207 162 209
rect 154 205 157 207
rect 159 205 162 207
rect 154 202 162 205
rect 164 210 172 212
rect 164 208 167 210
rect 169 208 172 210
rect 164 202 172 208
rect 174 208 179 215
rect 186 212 192 214
rect 186 210 188 212
rect 190 210 192 212
rect 186 208 192 210
rect 205 212 211 214
rect 205 210 207 212
rect 209 210 211 212
rect 205 208 211 210
rect 174 206 181 208
rect 174 204 177 206
rect 179 204 181 206
rect 174 202 181 204
rect 154 195 159 202
rect 186 201 191 208
rect 207 204 211 208
rect 207 201 213 204
rect 186 195 193 201
rect 195 199 203 201
rect 195 197 198 199
rect 200 197 203 199
rect 195 195 203 197
rect 205 195 213 201
rect 215 201 220 204
rect 215 199 222 201
rect 215 197 218 199
rect 220 197 222 199
rect 215 195 222 197
rect -71 96 -66 101
rect -73 94 -66 96
rect -73 92 -71 94
rect -69 92 -66 94
rect -73 90 -66 92
rect -64 90 -59 101
rect -57 92 -46 101
rect -44 98 -39 101
rect -44 96 -37 98
rect -31 96 -26 101
rect -44 94 -41 96
rect -39 94 -37 96
rect -44 92 -37 94
rect -33 94 -26 96
rect -33 92 -31 94
rect -29 92 -26 94
rect -57 90 -48 92
rect -55 84 -48 90
rect -33 90 -26 92
rect -24 90 -19 101
rect -17 92 -6 101
rect -4 98 1 101
rect -4 96 3 98
rect 29 96 34 103
rect -4 94 -1 96
rect 1 94 3 96
rect -4 92 3 94
rect 7 94 14 96
rect 7 92 9 94
rect 11 92 14 94
rect -17 90 -8 92
rect -55 82 -52 84
rect -50 82 -48 84
rect -55 80 -48 82
rect -15 84 -8 90
rect 7 90 14 92
rect -15 82 -12 84
rect -10 82 -8 84
rect -15 80 -8 82
rect 9 83 14 90
rect 16 90 24 96
rect 16 88 19 90
rect 21 88 24 90
rect 16 86 24 88
rect 26 93 34 96
rect 26 91 29 93
rect 31 91 34 93
rect 26 89 34 91
rect 36 101 44 103
rect 36 99 39 101
rect 41 99 44 101
rect 36 89 44 99
rect 46 101 53 103
rect 46 99 49 101
rect 51 99 53 101
rect 46 94 53 99
rect 59 96 64 103
rect 46 92 49 94
rect 51 92 53 94
rect 46 89 53 92
rect 57 94 64 96
rect 57 92 59 94
rect 61 92 64 94
rect 57 90 64 92
rect 26 86 31 89
rect 16 83 21 86
rect 59 83 64 90
rect 66 83 71 103
rect 73 97 80 103
rect 108 97 115 103
rect 73 87 82 97
rect 73 85 76 87
rect 78 85 82 87
rect 73 83 82 85
rect 84 94 91 97
rect 84 92 87 94
rect 89 92 91 94
rect 84 90 91 92
rect 97 94 104 97
rect 97 92 99 94
rect 101 92 104 94
rect 97 90 104 92
rect 84 83 89 90
rect 99 83 104 90
rect 106 87 115 97
rect 106 85 110 87
rect 112 85 115 87
rect 106 83 115 85
rect 117 83 122 103
rect 124 96 129 103
rect 135 101 142 103
rect 135 99 137 101
rect 139 99 142 101
rect 124 94 131 96
rect 124 92 127 94
rect 129 92 131 94
rect 124 90 131 92
rect 135 94 142 99
rect 135 92 137 94
rect 139 92 142 94
rect 124 83 129 90
rect 135 89 142 92
rect 144 101 152 103
rect 144 99 147 101
rect 149 99 152 101
rect 144 89 152 99
rect 154 96 159 103
rect 186 97 193 103
rect 195 101 203 103
rect 195 99 198 101
rect 200 99 203 101
rect 195 97 203 99
rect 205 97 213 103
rect 154 93 162 96
rect 154 91 157 93
rect 159 91 162 93
rect 154 89 162 91
rect 157 86 162 89
rect 164 90 172 96
rect 164 88 167 90
rect 169 88 172 90
rect 164 86 172 88
rect 167 83 172 86
rect 174 94 181 96
rect 174 92 177 94
rect 179 92 181 94
rect 174 90 181 92
rect 186 90 191 97
rect 207 94 213 97
rect 215 101 222 103
rect 215 99 218 101
rect 220 99 222 101
rect 215 97 222 99
rect 215 94 220 97
rect 207 90 211 94
rect 174 83 179 90
rect 186 88 192 90
rect 186 86 188 88
rect 190 86 192 88
rect 186 84 192 86
rect 205 88 211 90
rect 205 86 207 88
rect 209 86 211 88
rect 205 84 211 86
rect -55 72 -48 74
rect -55 70 -52 72
rect -50 70 -48 72
rect -55 64 -48 70
rect -15 72 -8 74
rect -15 70 -12 72
rect -10 70 -8 72
rect -73 62 -66 64
rect -73 60 -71 62
rect -69 60 -66 62
rect -73 58 -66 60
rect -71 53 -66 58
rect -64 53 -59 64
rect -57 62 -48 64
rect -15 64 -8 70
rect -33 62 -26 64
rect -57 53 -46 62
rect -44 60 -37 62
rect -44 58 -41 60
rect -39 58 -37 60
rect -33 60 -31 62
rect -29 60 -26 62
rect -33 58 -26 60
rect -44 56 -37 58
rect -44 53 -39 56
rect -31 53 -26 58
rect -24 53 -19 64
rect -17 62 -8 64
rect 9 64 14 71
rect 7 62 14 64
rect -17 53 -6 62
rect -4 60 3 62
rect -4 58 -1 60
rect 1 58 3 60
rect 7 60 9 62
rect 11 60 14 62
rect 7 58 14 60
rect 16 68 21 71
rect 16 66 24 68
rect 16 64 19 66
rect 21 64 24 66
rect 16 58 24 64
rect 26 65 31 68
rect 26 63 34 65
rect 26 61 29 63
rect 31 61 34 63
rect 26 58 34 61
rect -4 56 3 58
rect -4 53 1 56
rect 29 51 34 58
rect 36 55 44 65
rect 36 53 39 55
rect 41 53 44 55
rect 36 51 44 53
rect 46 62 53 65
rect 59 64 64 71
rect 46 60 49 62
rect 51 60 53 62
rect 46 55 53 60
rect 57 62 64 64
rect 57 60 59 62
rect 61 60 64 62
rect 57 58 64 60
rect 46 53 49 55
rect 51 53 53 55
rect 46 51 53 53
rect 59 51 64 58
rect 66 51 71 71
rect 73 69 82 71
rect 73 67 76 69
rect 78 67 82 69
rect 73 57 82 67
rect 84 64 89 71
rect 99 64 104 71
rect 84 62 91 64
rect 84 60 87 62
rect 89 60 91 62
rect 84 57 91 60
rect 97 62 104 64
rect 97 60 99 62
rect 101 60 104 62
rect 97 57 104 60
rect 106 69 115 71
rect 106 67 110 69
rect 112 67 115 69
rect 106 57 115 67
rect 73 51 80 57
rect 108 51 115 57
rect 117 51 122 71
rect 124 64 129 71
rect 167 68 172 71
rect 157 65 162 68
rect 124 62 131 64
rect 124 60 127 62
rect 129 60 131 62
rect 124 58 131 60
rect 135 62 142 65
rect 135 60 137 62
rect 139 60 142 62
rect 124 51 129 58
rect 135 55 142 60
rect 135 53 137 55
rect 139 53 142 55
rect 135 51 142 53
rect 144 55 152 65
rect 144 53 147 55
rect 149 53 152 55
rect 144 51 152 53
rect 154 63 162 65
rect 154 61 157 63
rect 159 61 162 63
rect 154 58 162 61
rect 164 66 172 68
rect 164 64 167 66
rect 169 64 172 66
rect 164 58 172 64
rect 174 64 179 71
rect 186 68 192 70
rect 186 66 188 68
rect 190 66 192 68
rect 186 64 192 66
rect 205 68 211 70
rect 205 66 207 68
rect 209 66 211 68
rect 205 64 211 66
rect 174 62 181 64
rect 174 60 177 62
rect 179 60 181 62
rect 174 58 181 60
rect 154 51 159 58
rect 186 57 191 64
rect 207 60 211 64
rect 207 57 213 60
rect 186 51 193 57
rect 195 55 203 57
rect 195 53 198 55
rect 200 53 203 55
rect 195 51 203 53
rect 205 51 213 57
rect 215 57 220 60
rect 215 55 222 57
rect 215 53 218 55
rect 220 53 222 55
rect 215 51 222 53
<< pdif >>
rect -73 278 -66 280
rect -73 276 -71 278
rect -69 276 -66 278
rect -73 267 -66 276
rect -64 278 -56 280
rect -64 276 -61 278
rect -59 276 -56 278
rect -64 271 -56 276
rect -64 269 -61 271
rect -59 269 -56 271
rect -64 267 -56 269
rect -54 278 -48 280
rect -33 278 -26 280
rect -54 276 -46 278
rect -54 274 -51 276
rect -49 274 -46 276
rect -54 267 -46 274
rect -52 260 -46 267
rect -44 273 -39 278
rect -33 276 -31 278
rect -29 276 -26 278
rect -44 271 -37 273
rect -44 269 -41 271
rect -39 269 -37 271
rect -44 264 -37 269
rect -33 267 -26 276
rect -24 278 -16 280
rect -24 276 -21 278
rect -19 276 -16 278
rect -24 271 -16 276
rect -24 269 -21 271
rect -19 269 -16 271
rect -24 267 -16 269
rect -14 278 -8 280
rect -14 276 -6 278
rect -14 274 -11 276
rect -9 274 -6 276
rect -14 267 -6 274
rect -44 262 -41 264
rect -39 262 -37 264
rect -44 260 -37 262
rect -12 260 -6 267
rect -4 273 1 278
rect 9 275 14 287
rect 7 273 14 275
rect -4 271 3 273
rect -4 269 -1 271
rect 1 269 3 271
rect -4 264 3 269
rect -4 262 -1 264
rect 1 262 3 264
rect 7 271 9 273
rect 11 271 14 273
rect 7 266 14 271
rect 7 264 9 266
rect 11 264 14 266
rect 7 262 14 264
rect 16 285 25 287
rect 16 283 20 285
rect 22 283 25 285
rect 48 285 62 287
rect 48 284 55 285
rect 16 275 25 283
rect 32 275 37 284
rect 16 262 27 275
rect 29 266 37 275
rect 29 264 32 266
rect 34 264 37 266
rect 29 262 37 264
rect -4 260 3 262
rect 32 259 37 262
rect 39 259 44 284
rect 46 283 55 284
rect 57 283 62 285
rect 46 278 62 283
rect 46 276 55 278
rect 57 276 62 278
rect 46 259 62 276
rect 64 277 72 287
rect 64 275 67 277
rect 69 275 72 277
rect 64 270 72 275
rect 64 268 67 270
rect 69 268 72 270
rect 64 259 72 268
rect 74 285 82 287
rect 74 283 77 285
rect 79 283 82 285
rect 74 278 82 283
rect 74 276 77 278
rect 79 276 82 278
rect 74 259 82 276
rect 84 272 89 287
rect 99 272 104 287
rect 84 270 91 272
rect 84 268 87 270
rect 89 268 91 270
rect 84 263 91 268
rect 84 261 87 263
rect 89 261 91 263
rect 84 259 91 261
rect 97 270 104 272
rect 97 268 99 270
rect 101 268 104 270
rect 97 263 104 268
rect 97 261 99 263
rect 101 261 104 263
rect 97 259 104 261
rect 106 285 114 287
rect 106 283 109 285
rect 111 283 114 285
rect 106 278 114 283
rect 106 276 109 278
rect 111 276 114 278
rect 106 259 114 276
rect 116 277 124 287
rect 116 275 119 277
rect 121 275 124 277
rect 116 270 124 275
rect 116 268 119 270
rect 121 268 124 270
rect 116 259 124 268
rect 126 285 140 287
rect 126 283 131 285
rect 133 284 140 285
rect 163 285 172 287
rect 133 283 142 284
rect 126 278 142 283
rect 126 276 131 278
rect 133 276 142 278
rect 126 259 142 276
rect 144 259 149 284
rect 151 275 156 284
rect 163 283 166 285
rect 168 283 172 285
rect 163 275 172 283
rect 151 266 159 275
rect 151 264 154 266
rect 156 264 159 266
rect 151 262 159 264
rect 161 262 172 275
rect 174 275 179 287
rect 188 280 193 287
rect 186 278 193 280
rect 186 276 188 278
rect 190 276 193 278
rect 174 273 181 275
rect 186 274 193 276
rect 174 271 177 273
rect 179 271 181 273
rect 174 266 181 271
rect 188 266 193 274
rect 195 266 200 287
rect 202 285 211 287
rect 202 283 207 285
rect 209 283 211 285
rect 202 277 211 283
rect 202 266 213 277
rect 174 264 177 266
rect 179 264 181 266
rect 174 262 181 264
rect 151 259 156 262
rect 205 259 213 266
rect 215 275 222 277
rect 215 273 218 275
rect 220 273 222 275
rect 215 268 222 273
rect 215 266 218 268
rect 220 266 222 268
rect 215 264 222 266
rect 215 259 220 264
rect -52 175 -46 182
rect -73 166 -66 175
rect -73 164 -71 166
rect -69 164 -66 166
rect -73 162 -66 164
rect -64 173 -56 175
rect -64 171 -61 173
rect -59 171 -56 173
rect -64 166 -56 171
rect -64 164 -61 166
rect -59 164 -56 166
rect -64 162 -56 164
rect -54 168 -46 175
rect -54 166 -51 168
rect -49 166 -46 168
rect -54 164 -46 166
rect -44 179 -37 182
rect -44 177 -41 179
rect -39 177 -37 179
rect -44 171 -37 177
rect -12 175 -6 182
rect -44 169 -41 171
rect -39 169 -37 171
rect -44 167 -37 169
rect -44 164 -39 167
rect -33 166 -26 175
rect -33 164 -31 166
rect -29 164 -26 166
rect -54 162 -48 164
rect -33 162 -26 164
rect -24 173 -16 175
rect -24 171 -21 173
rect -19 171 -16 173
rect -24 166 -16 171
rect -24 164 -21 166
rect -19 164 -16 166
rect -24 162 -16 164
rect -14 168 -6 175
rect -14 166 -11 168
rect -9 166 -6 168
rect -14 164 -6 166
rect -4 180 3 182
rect 32 180 37 183
rect -4 178 -1 180
rect 1 178 3 180
rect -4 173 3 178
rect -4 171 -1 173
rect 1 171 3 173
rect -4 169 3 171
rect 7 178 14 180
rect 7 176 9 178
rect 11 176 14 178
rect 7 171 14 176
rect 7 169 9 171
rect 11 169 14 171
rect -4 164 1 169
rect 7 167 14 169
rect -14 162 -8 164
rect 9 155 14 167
rect 16 167 27 180
rect 29 178 37 180
rect 29 176 32 178
rect 34 176 37 178
rect 29 167 37 176
rect 16 159 25 167
rect 16 157 20 159
rect 22 157 25 159
rect 32 158 37 167
rect 39 158 44 183
rect 46 166 62 183
rect 46 164 55 166
rect 57 164 62 166
rect 46 159 62 164
rect 46 158 55 159
rect 16 155 25 157
rect 48 157 55 158
rect 57 157 62 159
rect 48 155 62 157
rect 64 174 72 183
rect 64 172 67 174
rect 69 172 72 174
rect 64 167 72 172
rect 64 165 67 167
rect 69 165 72 167
rect 64 155 72 165
rect 74 166 82 183
rect 74 164 77 166
rect 79 164 82 166
rect 74 159 82 164
rect 74 157 77 159
rect 79 157 82 159
rect 74 155 82 157
rect 84 181 91 183
rect 84 179 87 181
rect 89 179 91 181
rect 84 174 91 179
rect 84 172 87 174
rect 89 172 91 174
rect 84 170 91 172
rect 97 181 104 183
rect 97 179 99 181
rect 101 179 104 181
rect 97 174 104 179
rect 97 172 99 174
rect 101 172 104 174
rect 97 170 104 172
rect 84 155 89 170
rect 99 155 104 170
rect 106 166 114 183
rect 106 164 109 166
rect 111 164 114 166
rect 106 159 114 164
rect 106 157 109 159
rect 111 157 114 159
rect 106 155 114 157
rect 116 174 124 183
rect 116 172 119 174
rect 121 172 124 174
rect 116 167 124 172
rect 116 165 119 167
rect 121 165 124 167
rect 116 155 124 165
rect 126 166 142 183
rect 126 164 131 166
rect 133 164 142 166
rect 126 159 142 164
rect 126 157 131 159
rect 133 158 142 159
rect 144 158 149 183
rect 151 180 156 183
rect 151 178 159 180
rect 151 176 154 178
rect 156 176 159 178
rect 151 167 159 176
rect 161 167 172 180
rect 151 158 156 167
rect 163 159 172 167
rect 133 157 140 158
rect 126 155 140 157
rect 163 157 166 159
rect 168 157 172 159
rect 163 155 172 157
rect 174 178 181 180
rect 174 176 177 178
rect 179 176 181 178
rect 205 176 213 183
rect 174 171 181 176
rect 174 169 177 171
rect 179 169 181 171
rect 174 167 181 169
rect 188 168 193 176
rect 174 155 179 167
rect 186 166 193 168
rect 186 164 188 166
rect 190 164 193 166
rect 186 162 193 164
rect 188 155 193 162
rect 195 155 200 176
rect 202 165 213 176
rect 215 178 220 183
rect 215 176 222 178
rect 215 174 218 176
rect 220 174 222 176
rect 215 169 222 174
rect 215 167 218 169
rect 220 167 222 169
rect 215 165 222 167
rect 202 159 211 165
rect 202 157 207 159
rect 209 157 211 159
rect 202 155 211 157
rect -73 134 -66 136
rect -73 132 -71 134
rect -69 132 -66 134
rect -73 123 -66 132
rect -64 134 -56 136
rect -64 132 -61 134
rect -59 132 -56 134
rect -64 127 -56 132
rect -64 125 -61 127
rect -59 125 -56 127
rect -64 123 -56 125
rect -54 134 -48 136
rect -33 134 -26 136
rect -54 132 -46 134
rect -54 130 -51 132
rect -49 130 -46 132
rect -54 123 -46 130
rect -52 116 -46 123
rect -44 132 -39 134
rect -33 132 -31 134
rect -29 132 -26 134
rect -44 130 -37 132
rect -44 128 -41 130
rect -39 128 -37 130
rect -44 122 -37 128
rect -33 123 -26 132
rect -24 134 -16 136
rect -24 132 -21 134
rect -19 132 -16 134
rect -24 127 -16 132
rect -24 125 -21 127
rect -19 125 -16 127
rect -24 123 -16 125
rect -14 134 -8 136
rect -14 132 -6 134
rect -14 130 -11 132
rect -9 130 -6 132
rect -14 123 -6 130
rect -44 120 -41 122
rect -39 120 -37 122
rect -44 116 -37 120
rect -12 116 -6 123
rect -4 129 1 134
rect 9 131 14 143
rect 7 129 14 131
rect -4 127 3 129
rect -4 125 -1 127
rect 1 125 3 127
rect -4 120 3 125
rect -4 118 -1 120
rect 1 118 3 120
rect 7 127 9 129
rect 11 127 14 129
rect 7 122 14 127
rect 7 120 9 122
rect 11 120 14 122
rect 7 118 14 120
rect 16 141 25 143
rect 16 139 20 141
rect 22 139 25 141
rect 48 141 62 143
rect 48 140 55 141
rect 16 131 25 139
rect 32 131 37 140
rect 16 118 27 131
rect 29 122 37 131
rect 29 120 32 122
rect 34 120 37 122
rect 29 118 37 120
rect -4 116 3 118
rect 32 115 37 118
rect 39 115 44 140
rect 46 139 55 140
rect 57 139 62 141
rect 46 134 62 139
rect 46 132 55 134
rect 57 132 62 134
rect 46 115 62 132
rect 64 133 72 143
rect 64 131 67 133
rect 69 131 72 133
rect 64 126 72 131
rect 64 124 67 126
rect 69 124 72 126
rect 64 115 72 124
rect 74 141 82 143
rect 74 139 77 141
rect 79 139 82 141
rect 74 134 82 139
rect 74 132 77 134
rect 79 132 82 134
rect 74 115 82 132
rect 84 128 89 143
rect 99 128 104 143
rect 84 126 91 128
rect 84 124 87 126
rect 89 124 91 126
rect 84 119 91 124
rect 84 117 87 119
rect 89 117 91 119
rect 84 115 91 117
rect 97 126 104 128
rect 97 124 99 126
rect 101 124 104 126
rect 97 119 104 124
rect 97 117 99 119
rect 101 117 104 119
rect 97 115 104 117
rect 106 141 114 143
rect 106 139 109 141
rect 111 139 114 141
rect 106 134 114 139
rect 106 132 109 134
rect 111 132 114 134
rect 106 115 114 132
rect 116 133 124 143
rect 116 131 119 133
rect 121 131 124 133
rect 116 126 124 131
rect 116 124 119 126
rect 121 124 124 126
rect 116 115 124 124
rect 126 141 140 143
rect 126 139 131 141
rect 133 140 140 141
rect 163 141 172 143
rect 133 139 142 140
rect 126 134 142 139
rect 126 132 131 134
rect 133 132 142 134
rect 126 115 142 132
rect 144 115 149 140
rect 151 131 156 140
rect 163 139 166 141
rect 168 139 172 141
rect 163 131 172 139
rect 151 122 159 131
rect 151 120 154 122
rect 156 120 159 122
rect 151 118 159 120
rect 161 118 172 131
rect 174 131 179 143
rect 188 136 193 143
rect 186 134 193 136
rect 186 132 188 134
rect 190 132 193 134
rect 174 129 181 131
rect 186 130 193 132
rect 174 127 177 129
rect 179 127 181 129
rect 174 122 181 127
rect 188 122 193 130
rect 195 122 200 143
rect 202 141 211 143
rect 202 139 207 141
rect 209 139 211 141
rect 202 133 211 139
rect 202 122 213 133
rect 174 120 177 122
rect 179 120 181 122
rect 174 118 181 120
rect 151 115 156 118
rect 205 115 213 122
rect 215 131 222 133
rect 215 129 218 131
rect 220 129 222 131
rect 215 124 222 129
rect 215 122 218 124
rect 220 122 222 124
rect 215 120 222 122
rect 215 115 220 120
rect -52 31 -46 38
rect -73 22 -66 31
rect -73 20 -71 22
rect -69 20 -66 22
rect -73 18 -66 20
rect -64 29 -56 31
rect -64 27 -61 29
rect -59 27 -56 29
rect -64 22 -56 27
rect -64 20 -61 22
rect -59 20 -56 22
rect -64 18 -56 20
rect -54 24 -46 31
rect -54 22 -51 24
rect -49 22 -46 24
rect -54 20 -46 22
rect -44 36 -37 38
rect -44 34 -41 36
rect -39 34 -37 36
rect -44 29 -37 34
rect -12 31 -6 38
rect -44 27 -41 29
rect -39 27 -37 29
rect -44 25 -37 27
rect -44 20 -39 25
rect -33 22 -26 31
rect -33 20 -31 22
rect -29 20 -26 22
rect -54 18 -48 20
rect -33 18 -26 20
rect -24 29 -16 31
rect -24 27 -21 29
rect -19 27 -16 29
rect -24 22 -16 27
rect -24 20 -21 22
rect -19 20 -16 22
rect -24 18 -16 20
rect -14 24 -6 31
rect -14 22 -11 24
rect -9 22 -6 24
rect -14 20 -6 22
rect -4 36 3 38
rect 32 36 37 39
rect -4 34 -1 36
rect 1 34 3 36
rect -4 29 3 34
rect -4 27 -1 29
rect 1 27 3 29
rect -4 25 3 27
rect 7 34 14 36
rect 7 32 9 34
rect 11 32 14 34
rect 7 27 14 32
rect 7 25 9 27
rect 11 25 14 27
rect -4 20 1 25
rect 7 23 14 25
rect -14 18 -8 20
rect 9 11 14 23
rect 16 23 27 36
rect 29 34 37 36
rect 29 32 32 34
rect 34 32 37 34
rect 29 23 37 32
rect 16 15 25 23
rect 16 13 20 15
rect 22 13 25 15
rect 32 14 37 23
rect 39 14 44 39
rect 46 22 62 39
rect 46 20 55 22
rect 57 20 62 22
rect 46 15 62 20
rect 46 14 55 15
rect 16 11 25 13
rect 48 13 55 14
rect 57 13 62 15
rect 48 11 62 13
rect 64 30 72 39
rect 64 28 67 30
rect 69 28 72 30
rect 64 23 72 28
rect 64 21 67 23
rect 69 21 72 23
rect 64 11 72 21
rect 74 22 82 39
rect 74 20 77 22
rect 79 20 82 22
rect 74 15 82 20
rect 74 13 77 15
rect 79 13 82 15
rect 74 11 82 13
rect 84 37 91 39
rect 84 35 87 37
rect 89 35 91 37
rect 84 30 91 35
rect 84 28 87 30
rect 89 28 91 30
rect 84 26 91 28
rect 97 37 104 39
rect 97 35 99 37
rect 101 35 104 37
rect 97 30 104 35
rect 97 28 99 30
rect 101 28 104 30
rect 97 26 104 28
rect 84 11 89 26
rect 99 11 104 26
rect 106 22 114 39
rect 106 20 109 22
rect 111 20 114 22
rect 106 15 114 20
rect 106 13 109 15
rect 111 13 114 15
rect 106 11 114 13
rect 116 30 124 39
rect 116 28 119 30
rect 121 28 124 30
rect 116 23 124 28
rect 116 21 119 23
rect 121 21 124 23
rect 116 11 124 21
rect 126 22 142 39
rect 126 20 131 22
rect 133 20 142 22
rect 126 15 142 20
rect 126 13 131 15
rect 133 14 142 15
rect 144 14 149 39
rect 151 36 156 39
rect 151 34 159 36
rect 151 32 154 34
rect 156 32 159 34
rect 151 23 159 32
rect 161 23 172 36
rect 151 14 156 23
rect 163 15 172 23
rect 133 13 140 14
rect 126 11 140 13
rect 163 13 166 15
rect 168 13 172 15
rect 163 11 172 13
rect 174 34 181 36
rect 174 32 177 34
rect 179 32 181 34
rect 205 32 213 39
rect 174 27 181 32
rect 174 25 177 27
rect 179 25 181 27
rect 174 23 181 25
rect 188 24 193 32
rect 174 11 179 23
rect 186 22 193 24
rect 186 20 188 22
rect 190 20 193 22
rect 186 18 193 20
rect 188 11 193 18
rect 195 11 200 32
rect 202 21 213 32
rect 215 34 220 39
rect 215 32 222 34
rect 215 30 218 32
rect 220 30 222 32
rect 215 25 222 30
rect 215 23 218 25
rect 220 23 222 25
rect 215 21 222 23
rect 202 15 211 21
rect 202 13 207 15
rect 209 13 211 15
rect 202 11 211 13
<< alu1 >>
rect -77 288 225 293
rect -77 286 -42 288
rect -40 286 -2 288
rect 0 286 217 288
rect 219 286 225 288
rect -77 285 225 286
rect -73 265 -69 272
rect -42 271 -37 273
rect -73 263 -72 265
rect -70 263 -69 265
rect -73 262 -60 263
rect -73 260 -68 262
rect -66 260 -60 262
rect -73 259 -60 260
rect -66 254 -52 255
rect -66 252 -58 254
rect -56 252 -52 254
rect -66 251 -52 252
rect -42 269 -41 271
rect -39 269 -37 271
rect -42 264 -37 269
rect -42 262 -41 264
rect -39 262 -37 264
rect -42 260 -37 262
rect -66 242 -61 251
rect -41 259 -37 260
rect -33 263 -29 272
rect 218 279 222 280
rect 209 275 222 279
rect 7 273 12 275
rect -2 271 3 273
rect -33 262 -20 263
rect -33 260 -28 262
rect -26 260 -20 262
rect -33 259 -20 260
rect -41 257 -40 259
rect -38 257 -37 259
rect -41 240 -37 257
rect -26 254 -12 255
rect -26 252 -18 254
rect -16 252 -12 254
rect -26 251 -12 252
rect -2 269 -1 271
rect 1 269 3 271
rect -2 264 3 269
rect -2 262 -1 264
rect 1 262 3 264
rect -2 260 3 262
rect -26 248 -21 251
rect -26 246 -24 248
rect -22 246 -21 248
rect -26 242 -21 246
rect -1 254 3 260
rect -1 252 0 254
rect 2 252 3 254
rect -49 238 -41 240
rect -39 238 -37 240
rect -1 240 3 252
rect -49 234 -37 238
rect -9 238 -1 240
rect 1 238 3 240
rect -9 234 3 238
rect 7 271 9 273
rect 11 271 12 273
rect 7 266 12 271
rect 7 264 9 266
rect 11 264 12 266
rect 7 262 12 264
rect 7 246 11 262
rect 38 262 76 263
rect 38 260 40 262
rect 42 260 76 262
rect 38 259 76 260
rect 38 256 43 259
rect 35 254 43 256
rect 35 252 36 254
rect 38 252 43 254
rect 35 250 43 252
rect 53 254 68 255
rect 53 252 55 254
rect 57 252 58 254
rect 60 252 62 254
rect 64 252 68 254
rect 53 251 68 252
rect 7 244 8 246
rect 10 244 11 246
rect 7 240 11 244
rect 7 238 12 240
rect 55 242 59 251
rect 86 270 92 272
rect 86 268 87 270
rect 89 268 92 270
rect 86 263 92 268
rect 86 261 87 263
rect 89 261 92 263
rect 86 259 92 261
rect 88 254 92 259
rect 88 252 89 254
rect 91 252 92 254
rect 88 239 92 252
rect 7 236 9 238
rect 11 236 12 238
rect 7 234 12 236
rect 86 238 92 239
rect 86 236 87 238
rect 89 236 92 238
rect 86 235 92 236
rect 96 270 102 272
rect 176 273 181 275
rect 176 271 177 273
rect 179 271 181 273
rect 96 268 99 270
rect 101 268 102 270
rect 96 267 102 268
rect 96 265 99 267
rect 101 265 102 267
rect 96 263 102 265
rect 96 261 99 263
rect 101 261 102 263
rect 96 259 102 261
rect 96 239 100 259
rect 112 262 150 263
rect 112 260 129 262
rect 131 260 150 262
rect 112 259 150 260
rect 145 256 150 259
rect 120 254 135 255
rect 120 252 124 254
rect 126 252 131 254
rect 133 252 135 254
rect 120 251 135 252
rect 145 254 153 256
rect 145 252 150 254
rect 152 252 153 254
rect 129 246 133 251
rect 145 250 153 252
rect 176 266 181 271
rect 176 264 177 266
rect 179 264 181 266
rect 176 262 181 264
rect 129 244 130 246
rect 132 244 133 246
rect 129 242 133 244
rect 96 238 102 239
rect 96 236 99 238
rect 101 236 102 238
rect 96 235 102 236
rect 177 240 181 262
rect 186 271 190 272
rect 186 269 187 271
rect 189 269 190 271
rect 186 263 190 269
rect 186 261 207 263
rect 186 259 191 261
rect 193 259 207 261
rect 186 254 207 255
rect 186 252 187 254
rect 189 252 201 254
rect 203 252 207 254
rect 186 251 207 252
rect 220 273 222 275
rect 218 268 222 273
rect 220 266 222 268
rect 186 242 190 251
rect 218 250 222 266
rect 218 248 219 250
rect 221 248 222 250
rect 218 247 222 248
rect 217 245 222 247
rect 217 243 218 245
rect 220 243 222 245
rect 217 241 222 243
rect 176 238 181 240
rect 176 236 177 238
rect 179 236 181 238
rect 176 234 181 236
rect -77 228 225 229
rect -77 226 -52 228
rect -50 226 -42 228
rect -40 226 -12 228
rect -10 226 -2 228
rect 0 226 217 228
rect 219 226 225 228
rect -77 225 225 226
rect -77 223 135 225
rect 137 223 225 225
rect -77 216 225 223
rect -77 214 -52 216
rect -50 214 -42 216
rect -40 214 -12 216
rect -10 214 -2 216
rect 0 214 217 216
rect 219 214 225 216
rect -77 213 225 214
rect -66 194 -61 200
rect -49 204 -37 208
rect -49 202 -41 204
rect -39 202 -37 204
rect -66 192 -64 194
rect -62 192 -61 194
rect -66 191 -61 192
rect -66 190 -52 191
rect -66 188 -58 190
rect -56 188 -52 190
rect -66 187 -52 188
rect -73 182 -60 183
rect -73 180 -68 182
rect -66 180 -60 182
rect -73 179 -60 180
rect -73 170 -69 179
rect -41 182 -37 202
rect -26 191 -21 200
rect -9 204 3 208
rect -9 202 -1 204
rect 1 202 3 204
rect -26 190 -12 191
rect -26 188 -18 190
rect -16 188 -12 190
rect -26 187 -12 188
rect -42 180 -40 182
rect -38 180 -37 182
rect -42 179 -37 180
rect -42 177 -41 179
rect -39 177 -37 179
rect -42 171 -37 177
rect -42 169 -41 171
rect -39 169 -37 171
rect -33 182 -20 183
rect -33 180 -28 182
rect -26 180 -20 182
rect -33 179 -20 180
rect -33 174 -29 179
rect -1 190 3 202
rect -1 188 0 190
rect 2 188 3 190
rect -1 182 3 188
rect -33 172 -32 174
rect -30 172 -29 174
rect -33 170 -29 172
rect -2 180 3 182
rect -2 178 -1 180
rect 1 178 3 180
rect -2 173 3 178
rect -42 167 -37 169
rect -2 171 -1 173
rect 1 171 3 173
rect -2 169 3 171
rect 7 206 12 208
rect 7 204 9 206
rect 11 204 12 206
rect 7 202 12 204
rect 7 198 11 202
rect 7 196 8 198
rect 10 196 11 198
rect 7 180 11 196
rect 86 206 92 207
rect 86 204 87 206
rect 89 204 92 206
rect 86 203 92 204
rect 7 178 12 180
rect 7 176 9 178
rect 11 176 12 178
rect 7 171 12 176
rect 35 190 43 192
rect 55 191 59 200
rect 35 188 36 190
rect 38 188 43 190
rect 35 186 43 188
rect 53 190 68 191
rect 53 188 55 190
rect 57 188 58 190
rect 60 188 62 190
rect 64 188 68 190
rect 53 187 68 188
rect 38 183 43 186
rect 88 190 92 203
rect 88 188 89 190
rect 91 188 92 190
rect 38 182 76 183
rect 38 180 53 182
rect 55 180 76 182
rect 38 179 76 180
rect 88 183 92 188
rect 86 181 92 183
rect 86 179 87 181
rect 89 179 92 181
rect 86 174 92 179
rect 86 172 87 174
rect 89 172 92 174
rect 7 169 9 171
rect 11 169 12 171
rect 7 167 12 169
rect 86 170 92 172
rect 96 206 102 207
rect 96 204 99 206
rect 101 204 102 206
rect 96 203 102 204
rect 176 206 183 208
rect 176 204 177 206
rect 179 204 183 206
rect 96 183 100 203
rect 129 198 133 200
rect 129 196 130 198
rect 132 196 133 198
rect 96 181 102 183
rect 96 179 99 181
rect 101 179 102 181
rect 96 177 102 179
rect 96 175 99 177
rect 101 175 102 177
rect 96 174 102 175
rect 96 172 99 174
rect 101 172 102 174
rect 96 170 102 172
rect 129 191 133 196
rect 176 202 183 204
rect 120 190 135 191
rect 120 188 124 190
rect 126 188 131 190
rect 133 188 135 190
rect 120 187 135 188
rect 145 190 153 192
rect 145 188 150 190
rect 152 188 153 190
rect 145 186 153 188
rect 145 185 150 186
rect 145 183 147 185
rect 149 183 150 185
rect 112 179 150 183
rect 177 180 181 202
rect 186 196 190 197
rect 186 194 187 196
rect 189 194 190 196
rect 186 191 190 194
rect 186 190 207 191
rect 186 188 201 190
rect 203 188 207 190
rect 186 187 207 188
rect 217 199 222 201
rect 217 197 218 199
rect 220 197 222 199
rect 217 195 222 197
rect 176 178 181 180
rect 176 176 177 178
rect 179 176 181 178
rect 176 171 181 176
rect 176 169 177 171
rect 179 169 181 171
rect 186 181 191 183
rect 193 181 207 183
rect 186 179 207 181
rect 186 177 190 179
rect 186 175 187 177
rect 189 175 190 177
rect 186 170 190 175
rect 176 167 181 169
rect 218 176 222 195
rect 220 174 222 176
rect 218 169 222 174
rect 220 167 222 169
rect 209 166 222 167
rect 209 164 211 166
rect 213 164 222 166
rect 209 163 222 164
rect 218 162 222 163
rect -77 156 225 157
rect -77 154 -42 156
rect -40 154 -2 156
rect 0 154 217 156
rect 219 154 225 156
rect -77 144 225 154
rect -77 142 -42 144
rect -40 142 -2 144
rect 0 142 217 144
rect 219 142 225 144
rect -77 141 225 142
rect -73 121 -69 128
rect -42 130 -37 132
rect -42 128 -41 130
rect -39 128 -37 130
rect -73 119 -72 121
rect -70 119 -69 121
rect -73 118 -60 119
rect -73 116 -68 118
rect -66 116 -60 118
rect -73 115 -60 116
rect -66 110 -52 111
rect -66 108 -58 110
rect -56 108 -52 110
rect -66 107 -52 108
rect -42 122 -37 128
rect -42 120 -41 122
rect -39 120 -37 122
rect -42 118 -37 120
rect -42 116 -40 118
rect -38 116 -37 118
rect -42 114 -37 116
rect -33 119 -29 128
rect 218 135 222 136
rect 209 131 222 135
rect 7 129 12 131
rect -2 127 3 129
rect -33 118 -20 119
rect -33 116 -28 118
rect -26 116 -20 118
rect -33 115 -20 116
rect -66 98 -61 107
rect -41 96 -37 114
rect -26 110 -12 111
rect -26 108 -18 110
rect -16 108 -12 110
rect -26 107 -12 108
rect -2 125 -1 127
rect 1 125 3 127
rect -2 120 3 125
rect -2 118 -1 120
rect 1 118 3 120
rect -2 116 3 118
rect -26 105 -21 107
rect -26 103 -24 105
rect -22 103 -21 105
rect -26 98 -21 103
rect -1 110 3 116
rect -1 108 0 110
rect 2 108 3 110
rect -49 94 -41 96
rect -39 94 -37 96
rect -1 96 3 108
rect -49 90 -37 94
rect -9 94 -1 96
rect 1 94 3 96
rect -9 90 3 94
rect 7 127 9 129
rect 11 127 12 129
rect 7 122 12 127
rect 7 120 9 122
rect 11 120 12 122
rect 7 118 12 120
rect 7 102 11 118
rect 38 118 76 119
rect 38 116 57 118
rect 59 116 76 118
rect 38 115 76 116
rect 38 112 43 115
rect 35 110 43 112
rect 35 108 36 110
rect 38 108 43 110
rect 35 106 43 108
rect 53 110 68 111
rect 53 108 55 110
rect 57 108 59 110
rect 61 108 62 110
rect 64 108 68 110
rect 53 107 68 108
rect 7 100 8 102
rect 10 100 11 102
rect 7 96 11 100
rect 7 94 12 96
rect 55 98 59 107
rect 86 126 92 128
rect 86 124 87 126
rect 89 124 92 126
rect 86 119 92 124
rect 86 117 87 119
rect 89 117 92 119
rect 86 115 92 117
rect 88 110 92 115
rect 88 108 89 110
rect 91 108 92 110
rect 88 95 92 108
rect 7 92 9 94
rect 11 92 12 94
rect 7 90 12 92
rect 86 94 92 95
rect 86 92 87 94
rect 89 92 92 94
rect 86 91 92 92
rect 96 126 102 128
rect 176 129 181 131
rect 176 127 177 129
rect 179 127 181 129
rect 96 124 99 126
rect 101 124 102 126
rect 96 123 102 124
rect 96 121 99 123
rect 101 121 102 123
rect 96 119 102 121
rect 96 117 99 119
rect 101 117 102 119
rect 96 115 102 117
rect 96 95 100 115
rect 112 118 150 119
rect 112 116 147 118
rect 149 116 150 118
rect 112 115 150 116
rect 145 112 150 115
rect 120 110 135 111
rect 120 108 124 110
rect 126 108 131 110
rect 133 108 135 110
rect 120 107 135 108
rect 145 110 153 112
rect 145 108 150 110
rect 152 108 153 110
rect 129 102 133 107
rect 145 106 153 108
rect 176 122 181 127
rect 176 120 177 122
rect 179 120 181 122
rect 176 118 181 120
rect 129 100 130 102
rect 132 100 133 102
rect 129 98 133 100
rect 96 94 102 95
rect 96 92 99 94
rect 101 92 102 94
rect 96 91 102 92
rect 177 96 181 118
rect 186 127 190 128
rect 186 125 187 127
rect 189 125 190 127
rect 186 119 190 125
rect 186 117 207 119
rect 186 115 191 117
rect 193 115 207 117
rect 186 110 207 111
rect 186 108 187 110
rect 189 108 201 110
rect 203 108 207 110
rect 186 107 207 108
rect 220 129 222 131
rect 218 124 222 129
rect 220 122 222 124
rect 186 103 190 107
rect 218 106 222 122
rect 218 104 219 106
rect 221 104 222 106
rect 218 103 222 104
rect 217 101 222 103
rect 217 99 218 101
rect 220 99 222 101
rect 217 97 222 99
rect 176 94 183 96
rect 176 92 177 94
rect 179 92 183 94
rect 176 90 183 92
rect -77 84 225 85
rect -77 82 -52 84
rect -50 82 -42 84
rect -40 82 -12 84
rect -10 82 -2 84
rect 0 82 217 84
rect 219 82 225 84
rect -77 75 225 82
rect -77 73 52 75
rect 54 73 225 75
rect -77 72 225 73
rect -77 70 -52 72
rect -50 70 -42 72
rect -40 70 -12 72
rect -10 70 -2 72
rect 0 70 217 72
rect 219 70 225 72
rect -77 69 225 70
rect -66 47 -61 56
rect -49 60 -37 64
rect -49 58 -41 60
rect -39 58 -37 60
rect -66 46 -52 47
rect -66 44 -58 46
rect -56 44 -52 46
rect -66 43 -52 44
rect -73 38 -60 39
rect -73 36 -68 38
rect -66 36 -60 38
rect -73 35 -60 36
rect -73 34 -69 35
rect -73 32 -72 34
rect -70 32 -69 34
rect -41 38 -37 58
rect -26 47 -21 56
rect -9 60 3 64
rect -9 58 -1 60
rect 1 58 3 60
rect -26 46 -12 47
rect -26 44 -18 46
rect -16 44 -12 46
rect -26 43 -12 44
rect -73 26 -69 32
rect -42 36 -37 38
rect -42 34 -41 36
rect -39 34 -37 36
rect -42 29 -37 34
rect -42 27 -41 29
rect -39 27 -37 29
rect -42 25 -37 27
rect -33 38 -20 39
rect -33 36 -28 38
rect -26 36 -20 38
rect -33 35 -20 36
rect -33 33 -29 35
rect -33 31 -32 33
rect -30 31 -29 33
rect -1 46 3 58
rect -1 44 0 46
rect 2 44 3 46
rect -1 38 3 44
rect -33 26 -29 31
rect -2 36 3 38
rect -2 34 -1 36
rect 1 34 3 36
rect -2 29 3 34
rect -2 27 -1 29
rect 1 27 3 29
rect -2 25 3 27
rect 7 62 12 64
rect 7 60 9 62
rect 11 60 12 62
rect 7 58 12 60
rect 7 54 11 58
rect 7 52 8 54
rect 10 52 11 54
rect 7 36 11 52
rect 86 62 92 63
rect 86 60 87 62
rect 89 60 92 62
rect 86 59 92 60
rect 7 34 12 36
rect 7 32 9 34
rect 11 32 12 34
rect 7 27 12 32
rect 35 46 43 48
rect 55 47 59 56
rect 35 44 36 46
rect 38 44 43 46
rect 35 42 43 44
rect 53 46 68 47
rect 53 44 55 46
rect 57 44 58 46
rect 60 44 62 46
rect 64 44 68 46
rect 53 43 68 44
rect 38 39 43 42
rect 88 46 92 59
rect 88 44 89 46
rect 91 44 92 46
rect 38 38 76 39
rect 38 36 52 38
rect 54 36 76 38
rect 38 35 76 36
rect 88 39 92 44
rect 86 37 92 39
rect 86 35 87 37
rect 89 35 92 37
rect 86 30 92 35
rect 86 28 87 30
rect 89 28 92 30
rect 7 25 9 27
rect 11 25 12 27
rect 7 23 12 25
rect 86 26 92 28
rect 96 62 102 63
rect 96 60 99 62
rect 101 60 102 62
rect 96 59 102 60
rect 176 62 183 64
rect 176 60 177 62
rect 179 60 183 62
rect 96 39 100 59
rect 129 54 133 56
rect 129 52 130 54
rect 132 52 133 54
rect 96 37 102 39
rect 96 35 99 37
rect 101 35 102 37
rect 96 33 102 35
rect 96 31 99 33
rect 101 31 102 33
rect 96 30 102 31
rect 96 28 99 30
rect 101 28 102 30
rect 96 26 102 28
rect 129 47 133 52
rect 176 58 183 60
rect 120 46 135 47
rect 120 44 124 46
rect 126 44 131 46
rect 133 44 135 46
rect 120 43 135 44
rect 145 46 153 48
rect 145 44 150 46
rect 152 44 153 46
rect 145 42 153 44
rect 145 41 150 42
rect 145 39 147 41
rect 149 39 150 41
rect 112 35 150 39
rect 177 36 181 58
rect 186 52 190 53
rect 186 50 187 52
rect 189 50 190 52
rect 186 47 190 50
rect 186 46 207 47
rect 186 44 201 46
rect 203 44 207 46
rect 186 43 207 44
rect 217 55 222 57
rect 217 53 218 55
rect 220 53 222 55
rect 217 51 222 53
rect 176 34 181 36
rect 176 32 177 34
rect 179 32 181 34
rect 176 27 181 32
rect 176 25 177 27
rect 179 25 181 27
rect 186 37 191 39
rect 193 37 207 39
rect 186 35 207 37
rect 186 33 190 35
rect 186 31 187 33
rect 189 31 190 33
rect 186 26 190 31
rect 176 23 181 25
rect 218 32 222 51
rect 220 30 222 32
rect 218 25 222 30
rect 220 23 222 25
rect 209 19 222 23
rect 218 18 222 19
rect -77 12 225 13
rect -77 10 -42 12
rect -40 10 -2 12
rect 0 10 217 12
rect 219 10 225 12
rect -77 5 225 10
<< alu2 >>
rect 102 271 190 272
rect 102 269 187 271
rect 189 269 190 271
rect 102 268 190 269
rect 98 267 106 268
rect -79 265 -69 266
rect -79 263 -78 265
rect -76 263 -72 265
rect -70 263 -69 265
rect 98 265 99 267
rect 101 265 106 267
rect 98 264 106 265
rect -79 262 -69 263
rect -36 262 43 263
rect -36 260 40 262
rect 42 260 43 262
rect -41 259 43 260
rect 128 262 136 263
rect 128 260 129 262
rect 131 260 132 262
rect 134 260 136 262
rect 128 259 136 260
rect -41 257 -40 259
rect -38 257 -32 259
rect -41 256 -32 257
rect -1 254 61 255
rect -1 252 0 254
rect 2 252 58 254
rect 60 252 61 254
rect -1 251 61 252
rect 88 254 191 255
rect 88 252 89 254
rect 91 252 187 254
rect 189 252 191 254
rect 88 251 191 252
rect 218 250 226 251
rect -37 248 -21 249
rect -37 246 -36 248
rect -34 246 -24 248
rect -22 246 -21 248
rect 218 248 219 250
rect 221 248 223 250
rect 225 248 226 250
rect 218 247 226 248
rect -37 244 -21 246
rect 7 246 133 247
rect 7 244 8 246
rect 10 244 130 246
rect 132 244 133 246
rect 7 243 133 244
rect 131 225 138 226
rect 131 223 132 225
rect 134 223 135 225
rect 137 223 138 225
rect 131 222 138 223
rect 7 198 133 199
rect 7 196 8 198
rect 10 196 130 198
rect 132 196 133 198
rect 7 195 133 196
rect 137 196 190 197
rect -79 194 -61 195
rect -79 192 -78 194
rect -76 192 -64 194
rect -62 192 -61 194
rect -79 191 -61 192
rect 137 194 187 196
rect 189 194 190 196
rect 137 193 190 194
rect 137 191 141 193
rect -1 190 61 191
rect -1 188 0 190
rect 2 188 58 190
rect 60 188 61 190
rect -1 187 61 188
rect 88 190 141 191
rect 88 188 89 190
rect 91 188 141 190
rect 88 187 141 188
rect 146 185 226 186
rect 146 183 147 185
rect 149 183 223 185
rect 225 183 226 185
rect -41 182 56 183
rect 146 182 226 183
rect -41 180 -40 182
rect -38 180 53 182
rect 55 180 56 182
rect -41 179 56 180
rect 98 177 190 178
rect 98 175 99 177
rect 101 175 187 177
rect 189 175 190 177
rect -37 174 -29 175
rect 98 174 190 175
rect -37 172 -36 174
rect -34 172 -32 174
rect -30 172 -29 174
rect -37 171 -29 172
rect 210 166 214 167
rect 210 164 211 166
rect 213 164 214 166
rect 138 127 190 128
rect 138 125 187 127
rect 189 125 190 127
rect 138 124 190 125
rect 98 123 142 124
rect -79 121 -69 122
rect -79 119 -78 121
rect -76 119 -72 121
rect -70 119 -69 121
rect 98 121 99 123
rect 101 121 142 123
rect 98 120 142 121
rect 210 119 214 164
rect -79 118 -69 119
rect -42 118 60 119
rect -42 116 -40 118
rect -38 116 57 118
rect 59 116 60 118
rect -42 115 60 116
rect 146 118 214 119
rect 146 116 147 118
rect 149 116 214 118
rect 146 115 214 116
rect -1 110 62 111
rect -1 108 0 110
rect 2 108 59 110
rect 61 108 62 110
rect -1 107 62 108
rect 88 110 191 111
rect 88 108 89 110
rect 91 108 187 110
rect 189 108 191 110
rect 88 107 191 108
rect 218 106 226 107
rect -37 105 -21 106
rect -37 103 -36 105
rect -34 103 -24 105
rect -22 103 -21 105
rect 218 104 219 106
rect 221 104 223 106
rect 225 104 226 106
rect 218 103 226 104
rect -37 102 -21 103
rect 7 102 133 103
rect 7 100 8 102
rect 10 100 130 102
rect 132 100 133 102
rect 7 99 133 100
rect 47 75 55 76
rect 47 73 48 75
rect 50 73 52 75
rect 54 73 55 75
rect 47 72 55 73
rect 7 54 133 55
rect 7 52 8 54
rect 10 52 130 54
rect 132 52 133 54
rect 7 51 133 52
rect 137 52 190 53
rect 137 50 187 52
rect 189 50 190 52
rect 137 49 190 50
rect 137 47 141 49
rect -1 46 61 47
rect -1 44 0 46
rect 2 44 58 46
rect 60 44 61 46
rect -1 43 61 44
rect 88 46 141 47
rect 88 44 89 46
rect 91 44 141 46
rect 88 43 141 44
rect 146 41 226 42
rect 146 39 147 41
rect 149 39 223 41
rect 225 39 226 41
rect 47 38 55 39
rect 146 38 226 39
rect 47 36 48 38
rect 50 36 52 38
rect 54 36 55 38
rect 47 35 55 36
rect -79 34 -69 35
rect -79 32 -78 34
rect -76 32 -72 34
rect -70 32 -69 34
rect -79 31 -69 32
rect -37 33 -29 34
rect -37 31 -36 33
rect -34 31 -32 33
rect -30 31 -29 33
rect -37 30 -29 31
rect 98 33 190 34
rect 98 31 99 33
rect 101 31 187 33
rect 189 31 190 33
rect 98 30 190 31
<< alu3 >>
rect -79 265 -75 266
rect -79 263 -78 265
rect -76 263 -75 265
rect -79 194 -75 263
rect 131 262 135 263
rect 131 260 132 262
rect 134 260 135 262
rect -79 192 -78 194
rect -76 192 -75 194
rect -79 121 -75 192
rect -79 119 -78 121
rect -76 119 -75 121
rect -79 34 -75 119
rect -79 32 -78 34
rect -76 32 -75 34
rect -79 28 -75 32
rect -37 248 -33 249
rect -37 246 -36 248
rect -34 246 -33 248
rect -37 174 -33 246
rect 131 225 135 260
rect 131 223 132 225
rect 134 223 135 225
rect 131 222 135 223
rect 222 250 226 251
rect 222 248 223 250
rect 225 248 226 250
rect 222 185 226 248
rect 222 183 223 185
rect 225 183 226 185
rect 222 182 226 183
rect -37 172 -36 174
rect -34 172 -33 174
rect -37 105 -33 172
rect -37 103 -36 105
rect -34 103 -33 105
rect -37 33 -33 103
rect 222 106 226 107
rect 222 104 223 106
rect 225 104 226 106
rect 47 75 51 76
rect 47 73 48 75
rect 50 73 51 75
rect 47 38 51 73
rect 222 41 226 104
rect 222 39 223 41
rect 225 39 226 41
rect 222 38 226 39
rect 47 36 48 38
rect 50 36 51 38
rect 47 35 51 36
rect -37 31 -36 33
rect -34 31 -33 33
rect -37 30 -33 31
<< ptie >>
rect -44 228 -38 230
rect -44 226 -42 228
rect -40 226 -38 228
rect -44 224 -38 226
rect -4 228 2 230
rect -4 226 -2 228
rect 0 226 2 228
rect -4 224 2 226
rect 215 228 221 230
rect 215 226 217 228
rect 219 226 221 228
rect 215 224 221 226
rect -44 216 -38 218
rect -44 214 -42 216
rect -40 214 -38 216
rect -44 212 -38 214
rect -4 216 2 218
rect -4 214 -2 216
rect 0 214 2 216
rect -4 212 2 214
rect 215 216 221 218
rect 215 214 217 216
rect 219 214 221 216
rect 215 212 221 214
rect -44 84 -38 86
rect -44 82 -42 84
rect -40 82 -38 84
rect -44 80 -38 82
rect -4 84 2 86
rect -4 82 -2 84
rect 0 82 2 84
rect -4 80 2 82
rect 215 84 221 86
rect 215 82 217 84
rect 219 82 221 84
rect 215 80 221 82
rect -44 72 -38 74
rect -44 70 -42 72
rect -40 70 -38 72
rect -44 68 -38 70
rect -4 72 2 74
rect -4 70 -2 72
rect 0 70 2 72
rect -4 68 2 70
rect 215 72 221 74
rect 215 70 217 72
rect 219 70 221 72
rect 215 68 221 70
<< ntie >>
rect -44 288 -38 290
rect -44 286 -42 288
rect -40 286 -38 288
rect -44 284 -38 286
rect -4 288 2 290
rect -4 286 -2 288
rect 0 286 2 288
rect -4 284 2 286
rect 215 288 221 290
rect 215 286 217 288
rect 219 286 221 288
rect 215 284 221 286
rect -44 156 -38 158
rect -44 154 -42 156
rect -40 154 -38 156
rect -44 152 -38 154
rect -4 156 2 158
rect -4 154 -2 156
rect 0 154 2 156
rect -4 152 2 154
rect 215 156 221 158
rect 215 154 217 156
rect 219 154 221 156
rect 215 152 221 154
rect -44 144 -38 146
rect -44 142 -42 144
rect -40 142 -38 144
rect -44 140 -38 142
rect -4 144 2 146
rect -4 142 -2 144
rect 0 142 2 144
rect -4 140 2 142
rect 215 144 221 146
rect 215 142 217 144
rect 219 142 221 144
rect 215 140 221 142
rect -44 12 -38 14
rect -44 10 -42 12
rect -40 10 -38 12
rect -44 8 -38 10
rect -4 12 2 14
rect -4 10 -2 12
rect 0 10 2 12
rect -4 8 2 10
rect 215 12 221 14
rect 215 10 217 12
rect 219 10 221 12
rect 215 8 221 10
<< nmos >>
rect -66 234 -64 245
rect -59 234 -57 245
rect -46 236 -44 245
rect -26 234 -24 245
rect -19 234 -17 245
rect -6 236 -4 245
rect 14 227 16 240
rect 24 230 26 240
rect 34 233 36 247
rect 44 233 46 247
rect 64 227 66 247
rect 71 227 73 247
rect 82 227 84 241
rect 104 227 106 241
rect 115 227 117 247
rect 122 227 124 247
rect 142 233 144 247
rect 152 233 154 247
rect 193 241 195 247
rect 203 241 205 247
rect 162 230 164 240
rect 172 227 174 240
rect 213 238 215 247
rect -66 197 -64 208
rect -59 197 -57 208
rect -46 197 -44 206
rect -26 197 -24 208
rect -19 197 -17 208
rect -6 197 -4 206
rect 14 202 16 215
rect 24 202 26 212
rect 34 195 36 209
rect 44 195 46 209
rect 64 195 66 215
rect 71 195 73 215
rect 82 201 84 215
rect 104 201 106 215
rect 115 195 117 215
rect 122 195 124 215
rect 142 195 144 209
rect 152 195 154 209
rect 162 202 164 212
rect 172 202 174 215
rect 193 195 195 201
rect 203 195 205 201
rect 213 195 215 204
rect -66 90 -64 101
rect -59 90 -57 101
rect -46 92 -44 101
rect -26 90 -24 101
rect -19 90 -17 101
rect -6 92 -4 101
rect 14 83 16 96
rect 24 86 26 96
rect 34 89 36 103
rect 44 89 46 103
rect 64 83 66 103
rect 71 83 73 103
rect 82 83 84 97
rect 104 83 106 97
rect 115 83 117 103
rect 122 83 124 103
rect 142 89 144 103
rect 152 89 154 103
rect 193 97 195 103
rect 203 97 205 103
rect 162 86 164 96
rect 172 83 174 96
rect 213 94 215 103
rect -66 53 -64 64
rect -59 53 -57 64
rect -46 53 -44 62
rect -26 53 -24 64
rect -19 53 -17 64
rect -6 53 -4 62
rect 14 58 16 71
rect 24 58 26 68
rect 34 51 36 65
rect 44 51 46 65
rect 64 51 66 71
rect 71 51 73 71
rect 82 57 84 71
rect 104 57 106 71
rect 115 51 117 71
rect 122 51 124 71
rect 142 51 144 65
rect 152 51 154 65
rect 162 58 164 68
rect 172 58 174 71
rect 193 51 195 57
rect 203 51 205 57
rect 213 51 215 60
<< pmos >>
rect -66 267 -64 280
rect -56 267 -54 280
rect -46 260 -44 278
rect -26 267 -24 280
rect -16 267 -14 280
rect -6 260 -4 278
rect 14 262 16 287
rect 27 262 29 275
rect 37 259 39 284
rect 44 259 46 284
rect 62 259 64 287
rect 72 259 74 287
rect 82 259 84 287
rect 104 259 106 287
rect 114 259 116 287
rect 124 259 126 287
rect 142 259 144 284
rect 149 259 151 284
rect 159 262 161 275
rect 172 262 174 287
rect 193 266 195 287
rect 200 266 202 287
rect 213 259 215 277
rect -66 162 -64 175
rect -56 162 -54 175
rect -46 164 -44 182
rect -26 162 -24 175
rect -16 162 -14 175
rect -6 164 -4 182
rect 14 155 16 180
rect 27 167 29 180
rect 37 158 39 183
rect 44 158 46 183
rect 62 155 64 183
rect 72 155 74 183
rect 82 155 84 183
rect 104 155 106 183
rect 114 155 116 183
rect 124 155 126 183
rect 142 158 144 183
rect 149 158 151 183
rect 159 167 161 180
rect 172 155 174 180
rect 193 155 195 176
rect 200 155 202 176
rect 213 165 215 183
rect -66 123 -64 136
rect -56 123 -54 136
rect -46 116 -44 134
rect -26 123 -24 136
rect -16 123 -14 136
rect -6 116 -4 134
rect 14 118 16 143
rect 27 118 29 131
rect 37 115 39 140
rect 44 115 46 140
rect 62 115 64 143
rect 72 115 74 143
rect 82 115 84 143
rect 104 115 106 143
rect 114 115 116 143
rect 124 115 126 143
rect 142 115 144 140
rect 149 115 151 140
rect 159 118 161 131
rect 172 118 174 143
rect 193 122 195 143
rect 200 122 202 143
rect 213 115 215 133
rect -66 18 -64 31
rect -56 18 -54 31
rect -46 20 -44 38
rect -26 18 -24 31
rect -16 18 -14 31
rect -6 20 -4 38
rect 14 11 16 36
rect 27 23 29 36
rect 37 14 39 39
rect 44 14 46 39
rect 62 11 64 39
rect 72 11 74 39
rect 82 11 84 39
rect 104 11 106 39
rect 114 11 116 39
rect 124 11 126 39
rect 142 14 144 39
rect 149 14 151 39
rect 159 23 161 36
rect 172 11 174 36
rect 193 11 195 32
rect 200 11 202 32
rect 213 21 215 39
<< polyct0 >>
rect -48 252 -46 254
rect -8 252 -6 254
rect 22 255 24 257
rect 16 245 18 247
rect 72 252 74 254
rect 82 252 84 254
rect 104 252 106 254
rect 114 252 116 254
rect 164 255 166 257
rect 211 252 213 254
rect 170 245 172 247
rect -48 188 -46 190
rect -8 188 -6 190
rect 16 195 18 197
rect 22 185 24 187
rect 72 188 74 190
rect 82 188 84 190
rect 104 188 106 190
rect 114 188 116 190
rect 170 195 172 197
rect 164 185 166 187
rect 211 188 213 190
rect -48 108 -46 110
rect -8 108 -6 110
rect 22 111 24 113
rect 16 101 18 103
rect 72 108 74 110
rect 82 108 84 110
rect 104 108 106 110
rect 114 108 116 110
rect 164 111 166 113
rect 211 108 213 110
rect 170 101 172 103
rect -48 44 -46 46
rect -8 44 -6 46
rect 16 51 18 53
rect 22 41 24 43
rect 72 44 74 46
rect 82 44 84 46
rect 104 44 106 46
rect 114 44 116 46
rect 170 51 172 53
rect 164 41 166 43
rect 211 44 213 46
<< polyct1 >>
rect -68 260 -66 262
rect -28 260 -26 262
rect -58 252 -56 254
rect -18 252 -16 254
rect 36 252 38 254
rect 55 252 57 254
rect 62 252 64 254
rect 124 252 126 254
rect 131 252 133 254
rect 150 252 152 254
rect 191 259 193 261
rect 201 252 203 254
rect -58 188 -56 190
rect -68 180 -66 182
rect -18 188 -16 190
rect -28 180 -26 182
rect 36 188 38 190
rect 55 188 57 190
rect 62 188 64 190
rect 124 188 126 190
rect 131 188 133 190
rect 150 188 152 190
rect 201 188 203 190
rect 191 181 193 183
rect -68 116 -66 118
rect -28 116 -26 118
rect -58 108 -56 110
rect -18 108 -16 110
rect 36 108 38 110
rect 55 108 57 110
rect 62 108 64 110
rect 124 108 126 110
rect 131 108 133 110
rect 150 108 152 110
rect 191 115 193 117
rect 201 108 203 110
rect -58 44 -56 46
rect -68 36 -66 38
rect -18 44 -16 46
rect -28 36 -26 38
rect 36 44 38 46
rect 55 44 57 46
rect 62 44 64 46
rect 124 44 126 46
rect 131 44 133 46
rect 150 44 152 46
rect 201 44 203 46
rect 191 37 193 39
<< ndifct0 >>
rect -71 236 -69 238
rect -31 236 -29 238
rect 19 232 21 234
rect 29 235 31 237
rect 39 243 41 245
rect 49 243 51 245
rect 49 236 51 238
rect 59 236 61 238
rect 76 229 78 231
rect 110 229 112 231
rect 137 243 139 245
rect 127 236 129 238
rect 137 236 139 238
rect 147 243 149 245
rect 198 243 200 245
rect 157 235 159 237
rect 167 232 169 234
rect 188 230 190 232
rect 207 230 209 232
rect -71 204 -69 206
rect -31 204 -29 206
rect 19 208 21 210
rect 29 205 31 207
rect 39 197 41 199
rect 49 204 51 206
rect 59 204 61 206
rect 49 197 51 199
rect 76 211 78 213
rect 110 211 112 213
rect 127 204 129 206
rect 137 204 139 206
rect 137 197 139 199
rect 147 197 149 199
rect 157 205 159 207
rect 167 208 169 210
rect 188 210 190 212
rect 207 210 209 212
rect 198 197 200 199
rect -71 92 -69 94
rect -31 92 -29 94
rect 19 88 21 90
rect 29 91 31 93
rect 39 99 41 101
rect 49 99 51 101
rect 49 92 51 94
rect 59 92 61 94
rect 76 85 78 87
rect 110 85 112 87
rect 137 99 139 101
rect 127 92 129 94
rect 137 92 139 94
rect 147 99 149 101
rect 198 99 200 101
rect 157 91 159 93
rect 167 88 169 90
rect 188 86 190 88
rect 207 86 209 88
rect -71 60 -69 62
rect -31 60 -29 62
rect 19 64 21 66
rect 29 61 31 63
rect 39 53 41 55
rect 49 60 51 62
rect 59 60 61 62
rect 49 53 51 55
rect 76 67 78 69
rect 110 67 112 69
rect 127 60 129 62
rect 137 60 139 62
rect 137 53 139 55
rect 147 53 149 55
rect 157 61 159 63
rect 167 64 169 66
rect 188 66 190 68
rect 207 66 209 68
rect 198 53 200 55
<< ndifct1 >>
rect -41 238 -39 240
rect -1 238 1 240
rect 9 236 11 238
rect -52 226 -50 228
rect -12 226 -10 228
rect 87 236 89 238
rect 99 236 101 238
rect 177 236 179 238
rect 218 243 220 245
rect -52 214 -50 216
rect -12 214 -10 216
rect -41 202 -39 204
rect -1 202 1 204
rect 9 204 11 206
rect 87 204 89 206
rect 99 204 101 206
rect 177 204 179 206
rect 218 197 220 199
rect -41 94 -39 96
rect -1 94 1 96
rect 9 92 11 94
rect -52 82 -50 84
rect -12 82 -10 84
rect 87 92 89 94
rect 99 92 101 94
rect 177 92 179 94
rect 218 99 220 101
rect -52 70 -50 72
rect -12 70 -10 72
rect -41 58 -39 60
rect -1 58 1 60
rect 9 60 11 62
rect 87 60 89 62
rect 99 60 101 62
rect 177 60 179 62
rect 218 53 220 55
<< ntiect1 >>
rect -42 286 -40 288
rect -2 286 0 288
rect 217 286 219 288
rect -42 154 -40 156
rect -2 154 0 156
rect 217 154 219 156
rect -42 142 -40 144
rect -2 142 0 144
rect 217 142 219 144
rect -42 10 -40 12
rect -2 10 0 12
rect 217 10 219 12
<< ptiect1 >>
rect -42 226 -40 228
rect -2 226 0 228
rect 217 226 219 228
rect -42 214 -40 216
rect -2 214 0 216
rect 217 214 219 216
rect -42 82 -40 84
rect -2 82 0 84
rect 217 82 219 84
rect -42 70 -40 72
rect -2 70 0 72
rect 217 70 219 72
<< pdifct0 >>
rect -71 276 -69 278
rect -61 276 -59 278
rect -61 269 -59 271
rect -51 274 -49 276
rect -31 276 -29 278
rect -21 276 -19 278
rect -21 269 -19 271
rect -11 274 -9 276
rect 20 283 22 285
rect 32 264 34 266
rect 55 283 57 285
rect 55 276 57 278
rect 67 275 69 277
rect 67 268 69 270
rect 77 283 79 285
rect 77 276 79 278
rect 109 283 111 285
rect 109 276 111 278
rect 119 275 121 277
rect 119 268 121 270
rect 131 283 133 285
rect 131 276 133 278
rect 166 283 168 285
rect 154 264 156 266
rect 188 276 190 278
rect 207 283 209 285
rect -71 164 -69 166
rect -61 171 -59 173
rect -61 164 -59 166
rect -51 166 -49 168
rect -31 164 -29 166
rect -21 171 -19 173
rect -21 164 -19 166
rect -11 166 -9 168
rect 32 176 34 178
rect 20 157 22 159
rect 55 164 57 166
rect 55 157 57 159
rect 67 172 69 174
rect 67 165 69 167
rect 77 164 79 166
rect 77 157 79 159
rect 109 164 111 166
rect 109 157 111 159
rect 119 172 121 174
rect 119 165 121 167
rect 131 164 133 166
rect 131 157 133 159
rect 154 176 156 178
rect 166 157 168 159
rect 188 164 190 166
rect 207 157 209 159
rect -71 132 -69 134
rect -61 132 -59 134
rect -61 125 -59 127
rect -51 130 -49 132
rect -31 132 -29 134
rect -21 132 -19 134
rect -21 125 -19 127
rect -11 130 -9 132
rect 20 139 22 141
rect 32 120 34 122
rect 55 139 57 141
rect 55 132 57 134
rect 67 131 69 133
rect 67 124 69 126
rect 77 139 79 141
rect 77 132 79 134
rect 109 139 111 141
rect 109 132 111 134
rect 119 131 121 133
rect 119 124 121 126
rect 131 139 133 141
rect 131 132 133 134
rect 166 139 168 141
rect 154 120 156 122
rect 188 132 190 134
rect 207 139 209 141
rect -71 20 -69 22
rect -61 27 -59 29
rect -61 20 -59 22
rect -51 22 -49 24
rect -31 20 -29 22
rect -21 27 -19 29
rect -21 20 -19 22
rect -11 22 -9 24
rect 32 32 34 34
rect 20 13 22 15
rect 55 20 57 22
rect 55 13 57 15
rect 67 28 69 30
rect 67 21 69 23
rect 77 20 79 22
rect 77 13 79 15
rect 109 20 111 22
rect 109 13 111 15
rect 119 28 121 30
rect 119 21 121 23
rect 131 20 133 22
rect 131 13 133 15
rect 154 32 156 34
rect 166 13 168 15
rect 188 20 190 22
rect 207 13 209 15
<< pdifct1 >>
rect -41 269 -39 271
rect -41 262 -39 264
rect -1 269 1 271
rect -1 262 1 264
rect 9 271 11 273
rect 9 264 11 266
rect 87 268 89 270
rect 87 261 89 263
rect 99 268 101 270
rect 99 261 101 263
rect 177 271 179 273
rect 177 264 179 266
rect 218 273 220 275
rect 218 266 220 268
rect -41 177 -39 179
rect -41 169 -39 171
rect -1 178 1 180
rect -1 171 1 173
rect 9 176 11 178
rect 9 169 11 171
rect 87 179 89 181
rect 87 172 89 174
rect 99 179 101 181
rect 99 172 101 174
rect 177 176 179 178
rect 177 169 179 171
rect 218 174 220 176
rect 218 167 220 169
rect -41 128 -39 130
rect -41 120 -39 122
rect -1 125 1 127
rect -1 118 1 120
rect 9 127 11 129
rect 9 120 11 122
rect 87 124 89 126
rect 87 117 89 119
rect 99 124 101 126
rect 99 117 101 119
rect 177 127 179 129
rect 177 120 179 122
rect 218 129 220 131
rect 218 122 220 124
rect -41 34 -39 36
rect -41 27 -39 29
rect -1 34 1 36
rect -1 27 1 29
rect 9 32 11 34
rect 9 25 11 27
rect 87 35 89 37
rect 87 28 89 30
rect 99 35 101 37
rect 99 28 101 30
rect 177 32 179 34
rect 177 25 179 27
rect 218 30 220 32
rect 218 23 220 25
<< alu0 >>
rect -73 278 -67 285
rect -73 276 -71 278
rect -69 276 -67 278
rect -73 275 -67 276
rect -62 278 -58 280
rect -62 276 -61 278
rect -59 276 -58 278
rect -62 271 -58 276
rect -53 276 -47 285
rect -53 274 -51 276
rect -49 274 -47 276
rect -33 278 -27 285
rect -33 276 -31 278
rect -29 276 -27 278
rect -33 275 -27 276
rect -22 278 -18 280
rect -22 276 -21 278
rect -19 276 -18 278
rect -53 273 -47 274
rect -62 269 -61 271
rect -59 270 -58 271
rect -59 269 -45 270
rect -62 266 -45 269
rect -49 254 -45 266
rect -49 252 -48 254
rect -46 252 -45 254
rect -49 247 -45 252
rect -57 243 -45 247
rect -22 271 -18 276
rect -13 276 -7 285
rect 18 283 20 285
rect 22 283 24 285
rect 18 282 24 283
rect 53 283 55 285
rect 57 283 59 285
rect -13 274 -11 276
rect -9 274 -7 276
rect 53 278 59 283
rect 75 283 77 285
rect 79 283 81 285
rect 53 276 55 278
rect 57 276 59 278
rect 53 275 59 276
rect 66 277 70 279
rect 66 275 67 277
rect 69 275 70 277
rect 75 278 81 283
rect 75 276 77 278
rect 79 276 81 278
rect 75 275 81 276
rect 107 283 109 285
rect 111 283 113 285
rect 107 278 113 283
rect 129 283 131 285
rect 133 283 135 285
rect 107 276 109 278
rect 111 276 113 278
rect 107 275 113 276
rect 118 277 122 279
rect 118 275 119 277
rect 121 275 122 277
rect 129 278 135 283
rect 164 283 166 285
rect 168 283 170 285
rect 164 282 170 283
rect 205 283 207 285
rect 209 283 211 285
rect 205 282 211 283
rect 129 276 131 278
rect 133 276 135 278
rect 129 275 135 276
rect 186 278 203 279
rect 186 276 188 278
rect 190 276 203 278
rect 186 275 203 276
rect -13 273 -7 274
rect -22 269 -21 271
rect -19 270 -18 271
rect -19 269 -5 270
rect -22 266 -5 269
rect -57 239 -53 243
rect -42 240 -41 242
rect -9 254 -5 266
rect -9 252 -8 254
rect -6 252 -5 254
rect -9 247 -5 252
rect -17 243 -5 247
rect -73 238 -53 239
rect -73 236 -71 238
rect -69 236 -53 238
rect -73 235 -53 236
rect -17 239 -13 243
rect -2 240 -1 242
rect -33 238 -13 239
rect -33 236 -31 238
rect -29 236 -13 238
rect -33 235 -13 236
rect 23 271 47 275
rect 66 271 70 275
rect 21 267 27 271
rect 43 270 83 271
rect 43 268 67 270
rect 69 268 83 270
rect 21 257 25 267
rect 31 266 35 268
rect 43 267 83 268
rect 31 264 32 266
rect 34 264 35 266
rect 31 263 35 264
rect 21 255 22 257
rect 24 255 25 257
rect 21 253 25 255
rect 28 259 35 263
rect 28 248 32 259
rect 71 254 75 259
rect 71 252 72 254
rect 74 252 75 254
rect 14 247 32 248
rect 14 245 16 247
rect 18 246 32 247
rect 18 245 43 246
rect 14 244 39 245
rect 28 243 39 244
rect 41 243 43 245
rect 28 242 43 243
rect 48 245 52 247
rect 48 243 49 245
rect 51 243 52 245
rect 48 238 52 243
rect 71 250 75 252
rect 79 256 83 267
rect 79 254 85 256
rect 79 252 82 254
rect 84 252 85 254
rect 79 250 85 252
rect 79 247 83 250
rect 63 243 83 247
rect 63 239 67 243
rect 27 237 49 238
rect 18 234 22 236
rect 27 235 29 237
rect 31 236 49 237
rect 51 236 52 238
rect 31 235 52 236
rect 57 238 67 239
rect 57 236 59 238
rect 61 236 67 238
rect 57 235 67 236
rect 118 271 122 275
rect 141 271 165 275
rect 105 270 145 271
rect 105 268 119 270
rect 121 268 145 270
rect 105 267 145 268
rect 105 256 109 267
rect 153 266 157 268
rect 161 267 167 271
rect 153 264 154 266
rect 156 264 157 266
rect 153 263 157 264
rect 153 259 160 263
rect 103 254 109 256
rect 103 252 104 254
rect 106 252 109 254
rect 103 250 109 252
rect 113 254 117 259
rect 113 252 114 254
rect 116 252 117 254
rect 113 250 117 252
rect 105 247 109 250
rect 105 243 125 247
rect 121 239 125 243
rect 156 248 160 259
rect 163 257 167 267
rect 163 255 164 257
rect 166 255 167 257
rect 163 253 167 255
rect 156 247 174 248
rect 136 245 140 247
rect 156 246 170 247
rect 136 243 137 245
rect 139 243 140 245
rect 121 238 131 239
rect 121 236 127 238
rect 129 236 131 238
rect 121 235 131 236
rect 136 238 140 243
rect 145 245 170 246
rect 172 245 174 247
rect 145 243 147 245
rect 149 244 174 245
rect 149 243 160 244
rect 145 242 160 243
rect 199 271 203 275
rect 199 267 214 271
rect 189 258 195 259
rect 210 254 214 267
rect 217 264 218 275
rect 210 252 211 254
rect 213 252 214 254
rect 210 246 214 252
rect 196 245 214 246
rect 196 243 198 245
rect 200 243 214 245
rect 196 242 214 243
rect 136 236 137 238
rect 139 237 161 238
rect 139 236 157 237
rect 136 235 157 236
rect 159 235 161 237
rect 27 234 52 235
rect 136 234 161 235
rect 166 234 170 236
rect 18 232 19 234
rect 21 232 22 234
rect 166 232 167 234
rect 169 232 170 234
rect 18 229 22 232
rect 74 231 80 232
rect 74 229 76 231
rect 78 229 80 231
rect 108 231 114 232
rect 108 229 110 231
rect 112 229 114 231
rect 166 229 170 232
rect 186 232 192 233
rect 186 230 188 232
rect 190 230 192 232
rect 186 229 192 230
rect 205 232 211 233
rect 205 230 207 232
rect 209 230 211 232
rect 205 229 211 230
rect 18 210 22 213
rect 74 211 76 213
rect 78 211 80 213
rect 74 210 80 211
rect 108 211 110 213
rect 112 211 114 213
rect 108 210 114 211
rect 166 210 170 213
rect 18 208 19 210
rect 21 208 22 210
rect 166 208 167 210
rect 169 208 170 210
rect 186 212 192 213
rect 186 210 188 212
rect 190 210 192 212
rect 186 209 192 210
rect 205 212 211 213
rect 205 210 207 212
rect 209 210 211 212
rect 205 209 211 210
rect -73 206 -53 207
rect -73 204 -71 206
rect -69 204 -53 206
rect -73 203 -53 204
rect -57 199 -53 203
rect -33 206 -13 207
rect -33 204 -31 206
rect -29 204 -13 206
rect -33 203 -13 204
rect -42 200 -41 202
rect -57 195 -45 199
rect -49 190 -45 195
rect -49 188 -48 190
rect -46 188 -45 190
rect -49 176 -45 188
rect -17 199 -13 203
rect -2 200 -1 202
rect -17 195 -5 199
rect -9 190 -5 195
rect -9 188 -8 190
rect -6 188 -5 190
rect -62 173 -45 176
rect -62 171 -61 173
rect -59 172 -45 173
rect -59 171 -58 172
rect -73 166 -67 167
rect -73 164 -71 166
rect -69 164 -67 166
rect -73 157 -67 164
rect -62 166 -58 171
rect -9 176 -5 188
rect -22 173 -5 176
rect -22 171 -21 173
rect -19 172 -5 173
rect -19 171 -18 172
rect -62 164 -61 166
rect -59 164 -58 166
rect -62 162 -58 164
rect -53 168 -47 169
rect -53 166 -51 168
rect -49 166 -47 168
rect -53 157 -47 166
rect -33 166 -27 167
rect -33 164 -31 166
rect -29 164 -27 166
rect -33 157 -27 164
rect -22 166 -18 171
rect 18 206 22 208
rect 27 207 52 208
rect 136 207 161 208
rect 27 205 29 207
rect 31 206 52 207
rect 31 205 49 206
rect 27 204 49 205
rect 51 204 52 206
rect 28 199 43 200
rect 28 198 39 199
rect 14 197 39 198
rect 41 197 43 199
rect 14 195 16 197
rect 18 196 43 197
rect 48 199 52 204
rect 57 206 67 207
rect 57 204 59 206
rect 61 204 67 206
rect 57 203 67 204
rect 48 197 49 199
rect 51 197 52 199
rect 18 195 32 196
rect 48 195 52 197
rect 14 194 32 195
rect 21 187 25 189
rect 21 185 22 187
rect 24 185 25 187
rect 21 175 25 185
rect 28 183 32 194
rect 63 199 67 203
rect 63 195 83 199
rect 79 192 83 195
rect 71 190 75 192
rect 71 188 72 190
rect 74 188 75 190
rect 71 183 75 188
rect 79 190 85 192
rect 79 188 82 190
rect 84 188 85 190
rect 79 186 85 188
rect 28 179 35 183
rect 31 178 35 179
rect 31 176 32 178
rect 34 176 35 178
rect 21 171 27 175
rect 31 174 35 176
rect 79 175 83 186
rect 43 174 83 175
rect 43 172 67 174
rect 69 172 83 174
rect 43 171 83 172
rect -22 164 -21 166
rect -19 164 -18 166
rect -22 162 -18 164
rect -13 168 -7 169
rect -13 166 -11 168
rect -9 166 -7 168
rect 23 167 47 171
rect 66 167 70 171
rect 121 206 131 207
rect 121 204 127 206
rect 129 204 131 206
rect 121 203 131 204
rect 136 206 157 207
rect 136 204 137 206
rect 139 205 157 206
rect 159 205 161 207
rect 166 206 170 208
rect 139 204 161 205
rect 121 199 125 203
rect 105 195 125 199
rect 105 192 109 195
rect 103 190 109 192
rect 103 188 104 190
rect 106 188 109 190
rect 103 186 109 188
rect 105 175 109 186
rect 113 190 117 192
rect 136 199 140 204
rect 136 197 137 199
rect 139 197 140 199
rect 136 195 140 197
rect 145 199 160 200
rect 145 197 147 199
rect 149 198 160 199
rect 149 197 174 198
rect 145 196 170 197
rect 156 195 170 196
rect 172 195 174 197
rect 156 194 174 195
rect 113 188 114 190
rect 116 188 117 190
rect 113 183 117 188
rect 156 183 160 194
rect 153 179 160 183
rect 163 187 167 189
rect 163 185 164 187
rect 166 185 167 187
rect 153 178 157 179
rect 153 176 154 178
rect 156 176 157 178
rect 105 174 145 175
rect 153 174 157 176
rect 163 175 167 185
rect 196 199 214 200
rect 196 197 198 199
rect 200 197 214 199
rect 196 196 214 197
rect 210 190 214 196
rect 210 188 211 190
rect 213 188 214 190
rect 189 183 195 184
rect 105 172 119 174
rect 121 172 145 174
rect 105 171 145 172
rect 161 171 167 175
rect 118 167 122 171
rect 141 167 165 171
rect 210 175 214 188
rect 199 171 214 175
rect 199 167 203 171
rect 217 167 218 178
rect -13 157 -7 166
rect 53 166 59 167
rect 53 164 55 166
rect 57 164 59 166
rect 18 159 24 160
rect 18 157 20 159
rect 22 157 24 159
rect 53 159 59 164
rect 66 165 67 167
rect 69 165 70 167
rect 66 163 70 165
rect 75 166 81 167
rect 75 164 77 166
rect 79 164 81 166
rect 53 157 55 159
rect 57 157 59 159
rect 75 159 81 164
rect 75 157 77 159
rect 79 157 81 159
rect 107 166 113 167
rect 107 164 109 166
rect 111 164 113 166
rect 107 159 113 164
rect 118 165 119 167
rect 121 165 122 167
rect 118 163 122 165
rect 129 166 135 167
rect 129 164 131 166
rect 133 164 135 166
rect 107 157 109 159
rect 111 157 113 159
rect 129 159 135 164
rect 186 166 203 167
rect 186 164 188 166
rect 190 164 203 166
rect 186 163 203 164
rect 129 157 131 159
rect 133 157 135 159
rect 164 159 170 160
rect 164 157 166 159
rect 168 157 170 159
rect 205 159 211 160
rect 205 157 207 159
rect 209 157 211 159
rect -73 134 -67 141
rect -73 132 -71 134
rect -69 132 -67 134
rect -73 131 -67 132
rect -62 134 -58 136
rect -62 132 -61 134
rect -59 132 -58 134
rect -62 127 -58 132
rect -53 132 -47 141
rect -33 134 -27 141
rect -33 132 -31 134
rect -29 132 -27 134
rect -53 130 -51 132
rect -49 130 -47 132
rect -53 129 -47 130
rect -33 131 -27 132
rect -22 134 -18 136
rect -22 132 -21 134
rect -19 132 -18 134
rect -62 125 -61 127
rect -59 126 -58 127
rect -59 125 -45 126
rect -62 122 -45 125
rect -49 110 -45 122
rect -22 127 -18 132
rect -13 132 -7 141
rect 18 139 20 141
rect 22 139 24 141
rect 18 138 24 139
rect 53 139 55 141
rect 57 139 59 141
rect -13 130 -11 132
rect -9 130 -7 132
rect 53 134 59 139
rect 75 139 77 141
rect 79 139 81 141
rect 53 132 55 134
rect 57 132 59 134
rect 53 131 59 132
rect 66 133 70 135
rect 66 131 67 133
rect 69 131 70 133
rect 75 134 81 139
rect 75 132 77 134
rect 79 132 81 134
rect 75 131 81 132
rect 107 139 109 141
rect 111 139 113 141
rect 107 134 113 139
rect 129 139 131 141
rect 133 139 135 141
rect 107 132 109 134
rect 111 132 113 134
rect 107 131 113 132
rect 118 133 122 135
rect 118 131 119 133
rect 121 131 122 133
rect 129 134 135 139
rect 164 139 166 141
rect 168 139 170 141
rect 164 138 170 139
rect 205 139 207 141
rect 209 139 211 141
rect 205 138 211 139
rect 129 132 131 134
rect 133 132 135 134
rect 129 131 135 132
rect 186 134 203 135
rect 186 132 188 134
rect 190 132 203 134
rect 186 131 203 132
rect -13 129 -7 130
rect -22 125 -21 127
rect -19 126 -18 127
rect -19 125 -5 126
rect -22 122 -5 125
rect -49 108 -48 110
rect -46 108 -45 110
rect -49 103 -45 108
rect -57 99 -45 103
rect -57 95 -53 99
rect -42 96 -41 98
rect -9 110 -5 122
rect -9 108 -8 110
rect -6 108 -5 110
rect -9 103 -5 108
rect -17 99 -5 103
rect -73 94 -53 95
rect -73 92 -71 94
rect -69 92 -53 94
rect -73 91 -53 92
rect -17 95 -13 99
rect -2 96 -1 98
rect -33 94 -13 95
rect -33 92 -31 94
rect -29 92 -13 94
rect -33 91 -13 92
rect 23 127 47 131
rect 66 127 70 131
rect 21 123 27 127
rect 43 126 83 127
rect 43 124 67 126
rect 69 124 83 126
rect 21 113 25 123
rect 31 122 35 124
rect 43 123 83 124
rect 31 120 32 122
rect 34 120 35 122
rect 31 119 35 120
rect 21 111 22 113
rect 24 111 25 113
rect 21 109 25 111
rect 28 115 35 119
rect 28 104 32 115
rect 71 110 75 115
rect 71 108 72 110
rect 74 108 75 110
rect 14 103 32 104
rect 14 101 16 103
rect 18 102 32 103
rect 18 101 43 102
rect 14 100 39 101
rect 28 99 39 100
rect 41 99 43 101
rect 28 98 43 99
rect 48 101 52 103
rect 48 99 49 101
rect 51 99 52 101
rect 48 94 52 99
rect 71 106 75 108
rect 79 112 83 123
rect 79 110 85 112
rect 79 108 82 110
rect 84 108 85 110
rect 79 106 85 108
rect 79 103 83 106
rect 63 99 83 103
rect 63 95 67 99
rect 27 93 49 94
rect 18 90 22 92
rect 27 91 29 93
rect 31 92 49 93
rect 51 92 52 94
rect 31 91 52 92
rect 57 94 67 95
rect 57 92 59 94
rect 61 92 67 94
rect 57 91 67 92
rect 118 127 122 131
rect 141 127 165 131
rect 105 126 145 127
rect 105 124 119 126
rect 121 124 145 126
rect 105 123 145 124
rect 105 112 109 123
rect 153 122 157 124
rect 161 123 167 127
rect 153 120 154 122
rect 156 120 157 122
rect 153 119 157 120
rect 153 115 160 119
rect 103 110 109 112
rect 103 108 104 110
rect 106 108 109 110
rect 103 106 109 108
rect 113 110 117 115
rect 113 108 114 110
rect 116 108 117 110
rect 113 106 117 108
rect 105 103 109 106
rect 105 99 125 103
rect 121 95 125 99
rect 156 104 160 115
rect 163 113 167 123
rect 163 111 164 113
rect 166 111 167 113
rect 163 109 167 111
rect 156 103 174 104
rect 136 101 140 103
rect 156 102 170 103
rect 136 99 137 101
rect 139 99 140 101
rect 121 94 131 95
rect 121 92 127 94
rect 129 92 131 94
rect 121 91 131 92
rect 136 94 140 99
rect 145 101 170 102
rect 172 101 174 103
rect 145 99 147 101
rect 149 100 174 101
rect 149 99 160 100
rect 145 98 160 99
rect 199 127 203 131
rect 199 123 214 127
rect 189 114 195 115
rect 210 110 214 123
rect 217 120 218 131
rect 210 108 211 110
rect 213 108 214 110
rect 210 102 214 108
rect 196 101 214 102
rect 196 99 198 101
rect 200 99 214 101
rect 196 98 214 99
rect 136 92 137 94
rect 139 93 161 94
rect 139 92 157 93
rect 136 91 157 92
rect 159 91 161 93
rect 27 90 52 91
rect 136 90 161 91
rect 166 90 170 92
rect 18 88 19 90
rect 21 88 22 90
rect 166 88 167 90
rect 169 88 170 90
rect 18 85 22 88
rect 74 87 80 88
rect 74 85 76 87
rect 78 85 80 87
rect 108 87 114 88
rect 108 85 110 87
rect 112 85 114 87
rect 166 85 170 88
rect 186 88 192 89
rect 186 86 188 88
rect 190 86 192 88
rect 186 85 192 86
rect 205 88 211 89
rect 205 86 207 88
rect 209 86 211 88
rect 205 85 211 86
rect 18 66 22 69
rect 74 67 76 69
rect 78 67 80 69
rect 74 66 80 67
rect 108 67 110 69
rect 112 67 114 69
rect 108 66 114 67
rect 166 66 170 69
rect 18 64 19 66
rect 21 64 22 66
rect 166 64 167 66
rect 169 64 170 66
rect 186 68 192 69
rect 186 66 188 68
rect 190 66 192 68
rect 186 65 192 66
rect 205 68 211 69
rect 205 66 207 68
rect 209 66 211 68
rect 205 65 211 66
rect -73 62 -53 63
rect -73 60 -71 62
rect -69 60 -53 62
rect -73 59 -53 60
rect -57 55 -53 59
rect -33 62 -13 63
rect -33 60 -31 62
rect -29 60 -13 62
rect -33 59 -13 60
rect -42 56 -41 58
rect -57 51 -45 55
rect -49 46 -45 51
rect -49 44 -48 46
rect -46 44 -45 46
rect -49 32 -45 44
rect -17 55 -13 59
rect -2 56 -1 58
rect -17 51 -5 55
rect -9 46 -5 51
rect -9 44 -8 46
rect -6 44 -5 46
rect -62 29 -45 32
rect -62 27 -61 29
rect -59 28 -45 29
rect -59 27 -58 28
rect -73 22 -67 23
rect -73 20 -71 22
rect -69 20 -67 22
rect -73 13 -67 20
rect -62 22 -58 27
rect -9 32 -5 44
rect -22 29 -5 32
rect -22 27 -21 29
rect -19 28 -5 29
rect -19 27 -18 28
rect -62 20 -61 22
rect -59 20 -58 22
rect -62 18 -58 20
rect -53 24 -47 25
rect -53 22 -51 24
rect -49 22 -47 24
rect -53 13 -47 22
rect -33 22 -27 23
rect -33 20 -31 22
rect -29 20 -27 22
rect -33 13 -27 20
rect -22 22 -18 27
rect 18 62 22 64
rect 27 63 52 64
rect 136 63 161 64
rect 27 61 29 63
rect 31 62 52 63
rect 31 61 49 62
rect 27 60 49 61
rect 51 60 52 62
rect 28 55 43 56
rect 28 54 39 55
rect 14 53 39 54
rect 41 53 43 55
rect 14 51 16 53
rect 18 52 43 53
rect 48 55 52 60
rect 57 62 67 63
rect 57 60 59 62
rect 61 60 67 62
rect 57 59 67 60
rect 48 53 49 55
rect 51 53 52 55
rect 18 51 32 52
rect 48 51 52 53
rect 14 50 32 51
rect 21 43 25 45
rect 21 41 22 43
rect 24 41 25 43
rect 21 31 25 41
rect 28 39 32 50
rect 63 55 67 59
rect 63 51 83 55
rect 79 48 83 51
rect 71 46 75 48
rect 71 44 72 46
rect 74 44 75 46
rect 71 39 75 44
rect 79 46 85 48
rect 79 44 82 46
rect 84 44 85 46
rect 79 42 85 44
rect 28 35 35 39
rect 31 34 35 35
rect 31 32 32 34
rect 34 32 35 34
rect 21 27 27 31
rect 31 30 35 32
rect 79 31 83 42
rect 43 30 83 31
rect 43 28 67 30
rect 69 28 83 30
rect 43 27 83 28
rect -22 20 -21 22
rect -19 20 -18 22
rect -22 18 -18 20
rect -13 24 -7 25
rect -13 22 -11 24
rect -9 22 -7 24
rect 23 23 47 27
rect 66 23 70 27
rect 121 62 131 63
rect 121 60 127 62
rect 129 60 131 62
rect 121 59 131 60
rect 136 62 157 63
rect 136 60 137 62
rect 139 61 157 62
rect 159 61 161 63
rect 166 62 170 64
rect 139 60 161 61
rect 121 55 125 59
rect 105 51 125 55
rect 105 48 109 51
rect 103 46 109 48
rect 103 44 104 46
rect 106 44 109 46
rect 103 42 109 44
rect 105 31 109 42
rect 113 46 117 48
rect 136 55 140 60
rect 136 53 137 55
rect 139 53 140 55
rect 136 51 140 53
rect 145 55 160 56
rect 145 53 147 55
rect 149 54 160 55
rect 149 53 174 54
rect 145 52 170 53
rect 156 51 170 52
rect 172 51 174 53
rect 156 50 174 51
rect 113 44 114 46
rect 116 44 117 46
rect 113 39 117 44
rect 156 39 160 50
rect 153 35 160 39
rect 163 43 167 45
rect 163 41 164 43
rect 166 41 167 43
rect 153 34 157 35
rect 153 32 154 34
rect 156 32 157 34
rect 105 30 145 31
rect 153 30 157 32
rect 163 31 167 41
rect 196 55 214 56
rect 196 53 198 55
rect 200 53 214 55
rect 196 52 214 53
rect 210 46 214 52
rect 210 44 211 46
rect 213 44 214 46
rect 189 39 195 40
rect 105 28 119 30
rect 121 28 145 30
rect 105 27 145 28
rect 161 27 167 31
rect 118 23 122 27
rect 141 23 165 27
rect 210 31 214 44
rect 199 27 214 31
rect 199 23 203 27
rect 217 23 218 34
rect -13 13 -7 22
rect 53 22 59 23
rect 53 20 55 22
rect 57 20 59 22
rect 18 15 24 16
rect 18 13 20 15
rect 22 13 24 15
rect 53 15 59 20
rect 66 21 67 23
rect 69 21 70 23
rect 66 19 70 21
rect 75 22 81 23
rect 75 20 77 22
rect 79 20 81 22
rect 53 13 55 15
rect 57 13 59 15
rect 75 15 81 20
rect 75 13 77 15
rect 79 13 81 15
rect 107 22 113 23
rect 107 20 109 22
rect 111 20 113 22
rect 107 15 113 20
rect 118 21 119 23
rect 121 21 122 23
rect 118 19 122 21
rect 129 22 135 23
rect 129 20 131 22
rect 133 20 135 22
rect 107 13 109 15
rect 111 13 113 15
rect 129 15 135 20
rect 186 22 203 23
rect 186 20 188 22
rect 190 20 203 22
rect 186 19 203 20
rect 129 13 131 15
rect 133 13 135 15
rect 164 15 170 16
rect 164 13 166 15
rect 168 13 170 15
rect 205 15 211 16
rect 205 13 207 15
rect 209 13 211 15
<< via1 >>
rect -72 263 -70 265
rect -40 257 -38 259
rect -24 246 -22 248
rect 0 252 2 254
rect 40 260 42 262
rect 58 252 60 254
rect 8 244 10 246
rect 89 252 91 254
rect 99 265 101 267
rect 129 260 131 262
rect 130 244 132 246
rect 187 269 189 271
rect 187 252 189 254
rect 219 248 221 250
rect 135 223 137 225
rect -64 192 -62 194
rect -40 180 -38 182
rect 0 188 2 190
rect -32 172 -30 174
rect 8 196 10 198
rect 58 188 60 190
rect 89 188 91 190
rect 53 180 55 182
rect 130 196 132 198
rect 99 175 101 177
rect 147 183 149 185
rect 187 194 189 196
rect 187 175 189 177
rect 211 164 213 166
rect -72 119 -70 121
rect -40 116 -38 118
rect -24 103 -22 105
rect 0 108 2 110
rect 57 116 59 118
rect 59 108 61 110
rect 8 100 10 102
rect 89 108 91 110
rect 99 121 101 123
rect 147 116 149 118
rect 130 100 132 102
rect 187 125 189 127
rect 187 108 189 110
rect 219 104 221 106
rect 52 73 54 75
rect -72 32 -70 34
rect -32 31 -30 33
rect 0 44 2 46
rect 8 52 10 54
rect 58 44 60 46
rect 89 44 91 46
rect 52 36 54 38
rect 130 52 132 54
rect 99 31 101 33
rect 147 39 149 41
rect 187 50 189 52
rect 187 31 189 33
<< via2 >>
rect -78 263 -76 265
rect 132 260 134 262
rect -36 246 -34 248
rect 223 248 225 250
rect 132 223 134 225
rect -78 192 -76 194
rect 223 183 225 185
rect -36 172 -34 174
rect -78 119 -76 121
rect -36 103 -34 105
rect 223 104 225 106
rect 48 73 50 75
rect 223 39 225 41
rect 48 36 50 38
rect -78 32 -76 34
rect -36 31 -34 33
<< labels >>
rlabel alu1 135 225 135 225 1 gnd
rlabel alu1 135 217 135 217 5 gnd
rlabel alu1 53 217 53 217 5 gnd
rlabel alu1 179 189 179 189 1 s_1
rlabel alu1 158 289 158 289 1 Vdd
rlabel alu1 184 289 184 289 1 Vdd
rlabel alu1 94 289 94 289 1 Vdd
rlabel alu1 29 289 29 289 1 vdd
rlabel alu1 29 152 29 152 1 Vdd
rlabel alu1 94 153 94 153 1 Vdd
rlabel alu1 185 153 185 153 1 Vdd
rlabel alu1 159 153 159 153 1 Vdd
rlabel alu1 159 9 159 9 1 Vdd
rlabel alu1 185 9 185 9 1 Vdd
rlabel alu1 94 9 94 9 1 Vdd
rlabel alu1 29 8 29 8 1 Vdd
rlabel alu1 29 145 29 145 1 vdd
rlabel alu1 94 145 94 145 1 Vdd
rlabel alu1 184 145 184 145 1 Vdd
rlabel alu1 158 145 158 145 1 Vdd
rlabel alu1 53 73 53 73 5 gnd
rlabel alu1 135 73 135 73 5 gnd
rlabel alu1 220 39 220 39 5 cout
rlabel alu1 135 81 135 81 1 gnd
rlabel alu1 53 81 53 81 1 gnd
rlabel alu1 179 114 179 114 1 s_2
rlabel alu1 179 45 179 45 1 s_3
rlabel alu1 -15 145 -15 145 4 vdd
rlabel alu1 -15 153 -15 153 2 vdd
rlabel alu1 -55 153 -55 153 2 vdd
rlabel alu1 -55 289 -55 289 4 vdd
rlabel alu1 -71 269 -71 269 1 b_0
rlabel alu1 -31 174 -31 174 1 b_1
rlabel alu1 -71 178 -71 178 1 a_2
rlabel via1 -63 193 -63 193 1 b_0
rlabel alu1 -63 247 -63 247 1 a_1
rlabel alu1 -23 193 -23 193 1 a_1
rlabel alu1 -55 145 -55 145 4 vdd
rlabel alu1 -71 121 -71 121 1 b_0
rlabel alu1 -63 104 -63 104 1 a_3
rlabel alu1 -23 105 -23 105 1 b_1
rlabel alu1 -31 121 -31 121 1 a_2
rlabel alu1 -71 32 -71 32 1 b_0
rlabel alu1 -63 49 -63 49 1 a_0
rlabel alu1 -39 44 -39 44 1 p_0
rlabel alu1 -23 49 -23 49 1 a_3
rlabel alu1 -31 33 -31 33 1 b_1
rlabel alu1 -31 265 -31 265 1 a_0
rlabel via1 -23 247 -23 247 1 b_1
rlabel alu1 179 258 179 258 1 p_1
<< end >>
