magic
tech scmos
timestamp 1519753522
<< nwell >>
rect -3465 133 -3453 148
<< polysilicon >>
rect -3460 141 -3458 143
rect -3460 131 -3458 138
rect -3459 127 -3458 131
rect -3460 122 -3458 127
rect -3460 117 -3458 119
<< ndiffusion >>
rect -3461 119 -3460 122
rect -3458 119 -3457 122
<< pdiffusion >>
rect -3461 138 -3460 141
rect -3458 138 -3457 141
<< metal1 >>
rect -3465 153 -3453 156
rect -3465 142 -3462 153
rect -3457 150 -3454 153
rect -3456 123 -3453 138
rect -3465 104 -3462 119
rect -3465 101 -3453 104
<< ntransistor >>
rect -3460 119 -3458 122
<< ptransistor >>
rect -3460 138 -3458 141
<< polycontact >>
rect -3463 127 -3459 131
<< ndcontact >>
rect -3465 119 -3461 123
rect -3457 119 -3453 123
<< pdcontact >>
rect -3465 138 -3461 142
rect -3457 138 -3453 142
<< nsubstratencontact >>
rect -3457 146 -3453 150
<< labels >>
rlabel metal1 -3460 155 -3460 155 5 vdd
rlabel metal1 -3460 102 -3460 102 1 gnd
rlabel polycontact -3461 129 -3461 129 3 in
rlabel metal1 -3454 129 -3454 129 7 out
<< end >>
