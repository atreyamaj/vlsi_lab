magic
tech scmos
timestamp 1555476560
<< nwell >>
rect -11 0 3 15
<< polysilicon >>
rect -5 7 -3 9
rect -5 -2 -3 1
rect -4 -6 -3 -2
rect -5 -9 -3 -6
rect -5 -14 -3 -12
<< ndiffusion >>
rect -6 -12 -5 -9
rect -3 -12 -2 -9
<< pdiffusion >>
rect -9 5 -5 7
rect -6 1 -5 5
rect -3 5 1 7
rect -3 1 -2 5
<< metal1 >>
rect -11 11 -1 15
rect -10 5 -6 11
rect -1 -9 2 1
rect -10 -17 -6 -13
rect -6 -21 2 -17
<< ntransistor >>
rect -5 -12 -3 -9
<< ptransistor >>
rect -5 1 -3 7
<< polycontact >>
rect -8 -6 -4 -2
<< ndcontact >>
rect -10 -13 -6 -9
rect -2 -13 2 -9
<< pdcontact >>
rect -10 1 -6 5
rect -2 1 2 5
<< psubstratepcontact >>
rect -10 -21 -6 -17
<< nsubstratencontact >>
rect -1 11 3 15
<< labels >>
rlabel metal1 1 -5 1 -5 7 out
rlabel polycontact -6 -4 -6 -4 1 in
rlabel metal1 -7 13 -7 13 4 Vdd
rlabel metal1 -3 -19 -3 -19 1 Gnd
<< end >>
