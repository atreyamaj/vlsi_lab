magic
tech scmos
timestamp 1553781431
<< ab >>
rect 5 63 134 77
rect 5 59 7 63
rect 9 59 134 63
rect 5 6 134 59
rect 5 -4 136 6
rect 5 -49 101 -4
rect 5 -53 97 -49
rect 99 -53 101 -49
rect 5 -67 101 -53
<< nwell >>
rect 0 37 139 82
rect 0 -72 106 -27
<< pwell >>
rect 0 0 139 37
rect 0 -4 136 0
rect 0 -27 106 -4
<< poly >>
rect 14 71 16 75
rect 37 68 39 73
rect 44 68 46 73
rect 62 71 64 75
rect 72 71 74 75
rect 82 71 84 75
rect 103 71 105 75
rect 110 71 112 75
rect 27 59 29 64
rect 14 33 16 46
rect 27 43 29 46
rect 123 61 125 66
rect 103 47 105 50
rect 99 45 105 47
rect 99 43 101 45
rect 103 43 105 45
rect 20 41 29 43
rect 20 39 22 41
rect 24 39 26 41
rect 37 40 39 43
rect 44 40 46 43
rect 62 40 64 43
rect 72 40 74 43
rect 82 40 84 43
rect 99 41 105 43
rect 20 37 26 39
rect 14 31 20 33
rect 14 29 16 31
rect 18 29 20 31
rect 14 27 20 29
rect 14 24 16 27
rect 24 24 26 37
rect 34 38 40 40
rect 34 36 36 38
rect 38 36 40 38
rect 34 34 40 36
rect 44 38 66 40
rect 44 36 55 38
rect 57 36 62 38
rect 64 36 66 38
rect 44 34 66 36
rect 70 38 76 40
rect 70 36 72 38
rect 74 36 76 38
rect 70 34 76 36
rect 80 38 86 40
rect 80 36 82 38
rect 84 36 86 38
rect 80 34 86 36
rect 34 31 36 34
rect 44 31 46 34
rect 64 31 66 34
rect 71 31 73 34
rect 14 7 16 11
rect 24 9 26 14
rect 34 12 36 17
rect 44 12 46 17
rect 82 25 84 34
rect 103 31 105 41
rect 110 40 112 50
rect 123 40 125 43
rect 109 38 115 40
rect 109 36 111 38
rect 113 36 115 38
rect 109 34 115 36
rect 119 38 125 40
rect 119 36 121 38
rect 123 36 125 38
rect 119 34 125 36
rect 113 31 115 34
rect 123 31 125 34
rect 103 20 105 25
rect 113 20 115 25
rect 123 17 125 22
rect 64 7 66 11
rect 71 7 73 11
rect 82 7 84 11
rect 22 -1 24 3
rect 33 -1 35 3
rect 40 -1 42 3
rect 22 -24 24 -15
rect 60 -7 62 -2
rect 70 -7 72 -2
rect 80 -4 82 1
rect 90 -1 92 3
rect 33 -24 35 -21
rect 40 -24 42 -21
rect 60 -24 62 -21
rect 70 -24 72 -21
rect 20 -26 26 -24
rect 20 -28 22 -26
rect 24 -28 26 -26
rect 20 -30 26 -28
rect 30 -26 36 -24
rect 30 -28 32 -26
rect 34 -28 36 -26
rect 30 -30 36 -28
rect 40 -26 62 -24
rect 40 -28 42 -26
rect 44 -28 49 -26
rect 51 -28 62 -26
rect 40 -30 62 -28
rect 66 -26 72 -24
rect 66 -28 68 -26
rect 70 -28 72 -26
rect 66 -30 72 -28
rect 80 -27 82 -14
rect 90 -17 92 -14
rect 86 -19 92 -17
rect 86 -21 88 -19
rect 90 -21 92 -19
rect 86 -23 92 -21
rect 80 -29 86 -27
rect 22 -33 24 -30
rect 32 -33 34 -30
rect 42 -33 44 -30
rect 60 -33 62 -30
rect 67 -33 69 -30
rect 80 -31 82 -29
rect 84 -31 86 -29
rect 77 -33 86 -31
rect 77 -36 79 -33
rect 90 -36 92 -23
rect 77 -54 79 -49
rect 22 -65 24 -61
rect 32 -65 34 -61
rect 42 -65 44 -61
rect 60 -63 62 -58
rect 67 -63 69 -58
rect 90 -65 92 -61
<< ndif >>
rect 29 24 34 31
rect 7 22 14 24
rect 7 20 9 22
rect 11 20 14 22
rect 7 18 14 20
rect 9 11 14 18
rect 16 18 24 24
rect 16 16 19 18
rect 21 16 24 18
rect 16 14 24 16
rect 26 21 34 24
rect 26 19 29 21
rect 31 19 34 21
rect 26 17 34 19
rect 36 29 44 31
rect 36 27 39 29
rect 41 27 44 29
rect 36 17 44 27
rect 46 29 53 31
rect 46 27 49 29
rect 51 27 53 29
rect 46 22 53 27
rect 59 24 64 31
rect 46 20 49 22
rect 51 20 53 22
rect 46 17 53 20
rect 57 22 64 24
rect 57 20 59 22
rect 61 20 64 22
rect 57 18 64 20
rect 26 14 31 17
rect 16 11 21 14
rect 59 11 64 18
rect 66 11 71 31
rect 73 25 80 31
rect 96 25 103 31
rect 105 29 113 31
rect 105 27 108 29
rect 110 27 113 29
rect 105 25 113 27
rect 115 25 123 31
rect 73 15 82 25
rect 73 13 76 15
rect 78 13 82 15
rect 73 11 82 13
rect 84 22 91 25
rect 84 20 87 22
rect 89 20 91 22
rect 84 18 91 20
rect 96 18 101 25
rect 117 22 123 25
rect 125 29 132 31
rect 125 27 128 29
rect 130 27 132 29
rect 125 25 132 27
rect 125 22 130 25
rect 117 18 121 22
rect 84 11 89 18
rect 96 16 102 18
rect 96 14 98 16
rect 100 14 102 16
rect 96 12 102 14
rect 115 16 121 18
rect 115 14 117 16
rect 119 14 121 16
rect 115 12 121 14
rect 17 -8 22 -1
rect 15 -10 22 -8
rect 15 -12 17 -10
rect 19 -12 22 -10
rect 15 -15 22 -12
rect 24 -3 33 -1
rect 24 -5 28 -3
rect 30 -5 33 -3
rect 24 -15 33 -5
rect 26 -21 33 -15
rect 35 -21 40 -1
rect 42 -8 47 -1
rect 85 -4 90 -1
rect 75 -7 80 -4
rect 42 -10 49 -8
rect 42 -12 45 -10
rect 47 -12 49 -10
rect 42 -14 49 -12
rect 53 -10 60 -7
rect 53 -12 55 -10
rect 57 -12 60 -10
rect 42 -21 47 -14
rect 53 -17 60 -12
rect 53 -19 55 -17
rect 57 -19 60 -17
rect 53 -21 60 -19
rect 62 -17 70 -7
rect 62 -19 65 -17
rect 67 -19 70 -17
rect 62 -21 70 -19
rect 72 -9 80 -7
rect 72 -11 75 -9
rect 77 -11 80 -9
rect 72 -14 80 -11
rect 82 -6 90 -4
rect 82 -8 85 -6
rect 87 -8 90 -6
rect 82 -14 90 -8
rect 92 -8 97 -1
rect 92 -10 99 -8
rect 92 -12 95 -10
rect 97 -12 99 -10
rect 92 -14 99 -12
rect 72 -21 77 -14
<< pdif >>
rect 9 59 14 71
rect 7 57 14 59
rect 7 55 9 57
rect 11 55 14 57
rect 7 50 14 55
rect 7 48 9 50
rect 11 48 14 50
rect 7 46 14 48
rect 16 69 25 71
rect 16 67 20 69
rect 22 67 25 69
rect 48 69 62 71
rect 48 68 55 69
rect 16 59 25 67
rect 32 59 37 68
rect 16 46 27 59
rect 29 50 37 59
rect 29 48 32 50
rect 34 48 37 50
rect 29 46 37 48
rect 32 43 37 46
rect 39 43 44 68
rect 46 67 55 68
rect 57 67 62 69
rect 46 62 62 67
rect 46 60 55 62
rect 57 60 62 62
rect 46 43 62 60
rect 64 61 72 71
rect 64 59 67 61
rect 69 59 72 61
rect 64 54 72 59
rect 64 52 67 54
rect 69 52 72 54
rect 64 43 72 52
rect 74 69 82 71
rect 74 67 77 69
rect 79 67 82 69
rect 74 62 82 67
rect 74 60 77 62
rect 79 60 82 62
rect 74 43 82 60
rect 84 56 89 71
rect 98 64 103 71
rect 96 62 103 64
rect 96 60 98 62
rect 100 60 103 62
rect 96 58 103 60
rect 84 54 91 56
rect 84 52 87 54
rect 89 52 91 54
rect 84 47 91 52
rect 98 50 103 58
rect 105 50 110 71
rect 112 69 121 71
rect 112 67 117 69
rect 119 67 121 69
rect 112 61 121 67
rect 112 50 123 61
rect 84 45 87 47
rect 89 45 91 47
rect 84 43 91 45
rect 115 43 123 50
rect 125 59 132 61
rect 125 57 128 59
rect 130 57 132 59
rect 125 52 132 57
rect 125 50 128 52
rect 130 50 132 52
rect 125 48 132 50
rect 125 43 130 48
rect 15 -35 22 -33
rect 15 -37 17 -35
rect 19 -37 22 -35
rect 15 -42 22 -37
rect 15 -44 17 -42
rect 19 -44 22 -42
rect 15 -46 22 -44
rect 17 -61 22 -46
rect 24 -50 32 -33
rect 24 -52 27 -50
rect 29 -52 32 -50
rect 24 -57 32 -52
rect 24 -59 27 -57
rect 29 -59 32 -57
rect 24 -61 32 -59
rect 34 -42 42 -33
rect 34 -44 37 -42
rect 39 -44 42 -42
rect 34 -49 42 -44
rect 34 -51 37 -49
rect 39 -51 42 -49
rect 34 -61 42 -51
rect 44 -50 60 -33
rect 44 -52 49 -50
rect 51 -52 60 -50
rect 44 -57 60 -52
rect 44 -59 49 -57
rect 51 -58 60 -57
rect 62 -58 67 -33
rect 69 -36 74 -33
rect 69 -38 77 -36
rect 69 -40 72 -38
rect 74 -40 77 -38
rect 69 -49 77 -40
rect 79 -49 90 -36
rect 69 -58 74 -49
rect 81 -57 90 -49
rect 51 -59 58 -58
rect 44 -61 58 -59
rect 81 -59 84 -57
rect 86 -59 90 -57
rect 81 -61 90 -59
rect 92 -38 99 -36
rect 92 -40 95 -38
rect 97 -40 99 -38
rect 92 -45 99 -40
rect 92 -47 95 -45
rect 97 -47 99 -45
rect 92 -49 99 -47
rect 92 -61 97 -49
<< alu1 >>
rect 3 72 136 77
rect 3 70 127 72
rect 129 70 136 72
rect 3 69 136 70
rect 128 63 132 64
rect 119 59 132 63
rect 7 57 12 59
rect 7 55 9 57
rect 11 55 12 57
rect 7 50 12 55
rect 7 48 9 50
rect 11 48 12 50
rect 7 46 12 48
rect 7 33 11 46
rect 38 43 76 47
rect 7 31 8 33
rect 10 31 11 33
rect 38 40 43 43
rect 35 38 43 40
rect 35 36 36 38
rect 38 36 43 38
rect 35 34 43 36
rect 53 38 68 39
rect 53 36 55 38
rect 57 36 62 38
rect 64 36 68 38
rect 53 35 68 36
rect 7 24 11 31
rect 7 22 12 24
rect 55 26 59 35
rect 86 54 92 56
rect 86 52 87 54
rect 89 52 92 54
rect 96 52 100 56
rect 86 48 100 52
rect 86 47 92 48
rect 86 45 87 47
rect 89 45 92 47
rect 86 43 92 45
rect 96 47 100 48
rect 96 45 117 47
rect 96 43 101 45
rect 103 43 117 45
rect 88 23 92 43
rect 96 38 117 39
rect 96 36 111 38
rect 113 36 117 38
rect 96 35 117 36
rect 130 57 132 59
rect 128 52 132 57
rect 130 50 132 52
rect 96 33 100 35
rect 96 31 97 33
rect 99 31 100 33
rect 96 26 100 31
rect 128 31 132 50
rect 127 29 132 31
rect 127 27 128 29
rect 130 27 132 29
rect 127 25 132 27
rect 7 20 9 22
rect 11 20 12 22
rect 7 18 12 20
rect 86 22 92 23
rect 86 20 87 22
rect 89 20 92 22
rect 86 19 92 20
rect 3 12 136 13
rect 3 10 127 12
rect 129 10 136 12
rect 3 -3 136 10
rect 14 -10 20 -9
rect 14 -12 17 -10
rect 19 -12 20 -10
rect 14 -13 20 -12
rect 94 -10 99 -8
rect 94 -12 95 -10
rect 97 -12 99 -10
rect 14 -33 18 -13
rect 47 -20 51 -16
rect 47 -22 48 -20
rect 50 -22 51 -20
rect 94 -14 99 -12
rect 14 -35 20 -33
rect 14 -37 17 -35
rect 19 -37 20 -35
rect 14 -38 20 -37
rect 14 -40 17 -38
rect 19 -40 20 -38
rect 14 -42 20 -40
rect 14 -44 17 -42
rect 19 -44 20 -42
rect 14 -46 20 -44
rect 47 -25 51 -22
rect 38 -26 53 -25
rect 38 -28 42 -26
rect 44 -28 49 -26
rect 51 -28 53 -26
rect 38 -29 53 -28
rect 63 -26 71 -24
rect 63 -28 68 -26
rect 70 -28 71 -26
rect 63 -30 71 -28
rect 63 -33 68 -30
rect 30 -37 68 -33
rect 95 -36 99 -14
rect 94 -38 99 -36
rect 94 -40 95 -38
rect 97 -40 99 -38
rect 94 -45 99 -40
rect 94 -47 95 -45
rect 97 -47 99 -45
rect 94 -49 99 -47
rect 3 -67 103 -59
<< alu2 >>
rect 7 33 11 36
rect 7 31 8 33
rect 10 31 11 33
rect 7 -19 11 31
rect 96 33 100 34
rect 96 31 97 33
rect 99 31 100 33
rect 7 -20 51 -19
rect 7 -22 48 -20
rect 50 -22 51 -20
rect 7 -23 51 -22
rect 96 -37 100 31
rect 16 -38 100 -37
rect 16 -40 17 -38
rect 19 -40 100 -38
rect 16 -41 100 -40
<< ptie >>
rect 125 12 131 14
rect 125 10 127 12
rect 129 10 131 12
rect 125 8 131 10
<< ntie >>
rect 125 72 131 74
rect 125 70 127 72
rect 129 70 131 72
rect 125 68 131 70
<< nmos >>
rect 14 11 16 24
rect 24 14 26 24
rect 34 17 36 31
rect 44 17 46 31
rect 64 11 66 31
rect 71 11 73 31
rect 103 25 105 31
rect 113 25 115 31
rect 82 11 84 25
rect 123 22 125 31
rect 22 -15 24 -1
rect 33 -21 35 -1
rect 40 -21 42 -1
rect 60 -21 62 -7
rect 70 -21 72 -7
rect 80 -14 82 -4
rect 90 -14 92 -1
<< pmos >>
rect 14 46 16 71
rect 27 46 29 59
rect 37 43 39 68
rect 44 43 46 68
rect 62 43 64 71
rect 72 43 74 71
rect 82 43 84 71
rect 103 50 105 71
rect 110 50 112 71
rect 123 43 125 61
rect 22 -61 24 -33
rect 32 -61 34 -33
rect 42 -61 44 -33
rect 60 -58 62 -33
rect 67 -58 69 -33
rect 77 -49 79 -36
rect 90 -61 92 -36
<< polyct0 >>
rect 22 39 24 41
rect 16 29 18 31
rect 72 36 74 38
rect 82 36 84 38
rect 121 36 123 38
rect 22 -28 24 -26
rect 32 -28 34 -26
rect 88 -21 90 -19
rect 82 -31 84 -29
<< polyct1 >>
rect 101 43 103 45
rect 36 36 38 38
rect 55 36 57 38
rect 62 36 64 38
rect 111 36 113 38
rect 42 -28 44 -26
rect 49 -28 51 -26
rect 68 -28 70 -26
<< ndifct0 >>
rect 19 16 21 18
rect 29 19 31 21
rect 39 27 41 29
rect 49 27 51 29
rect 49 20 51 22
rect 59 20 61 22
rect 108 27 110 29
rect 76 13 78 15
rect 98 14 100 16
rect 117 14 119 16
rect 28 -5 30 -3
rect 45 -12 47 -10
rect 55 -12 57 -10
rect 55 -19 57 -17
rect 65 -19 67 -17
rect 75 -11 77 -9
rect 85 -8 87 -6
<< ndifct1 >>
rect 9 20 11 22
rect 87 20 89 22
rect 128 27 130 29
rect 17 -12 19 -10
rect 95 -12 97 -10
<< ntiect1 >>
rect 127 70 129 72
<< ptiect1 >>
rect 127 10 129 12
<< pdifct0 >>
rect 20 67 22 69
rect 32 48 34 50
rect 55 67 57 69
rect 55 60 57 62
rect 67 59 69 61
rect 67 52 69 54
rect 77 67 79 69
rect 77 60 79 62
rect 98 60 100 62
rect 117 67 119 69
rect 27 -52 29 -50
rect 27 -59 29 -57
rect 37 -44 39 -42
rect 37 -51 39 -49
rect 49 -52 51 -50
rect 49 -59 51 -57
rect 72 -40 74 -38
rect 84 -59 86 -57
<< pdifct1 >>
rect 9 55 11 57
rect 9 48 11 50
rect 87 52 89 54
rect 87 45 89 47
rect 128 57 130 59
rect 128 50 130 52
rect 17 -37 19 -35
rect 17 -44 19 -42
rect 95 -40 97 -38
rect 95 -47 97 -45
<< alu0 >>
rect 18 67 20 69
rect 22 67 24 69
rect 18 66 24 67
rect 53 67 55 69
rect 57 67 59 69
rect 53 62 59 67
rect 75 67 77 69
rect 79 67 81 69
rect 53 60 55 62
rect 57 60 59 62
rect 53 59 59 60
rect 66 61 70 63
rect 66 59 67 61
rect 69 59 70 61
rect 75 62 81 67
rect 115 67 117 69
rect 119 67 121 69
rect 115 66 121 67
rect 75 60 77 62
rect 79 60 81 62
rect 75 59 81 60
rect 96 62 113 63
rect 96 60 98 62
rect 100 60 113 62
rect 96 59 113 60
rect 23 55 47 59
rect 66 55 70 59
rect 21 51 27 55
rect 43 54 83 55
rect 43 52 67 54
rect 69 52 83 54
rect 21 41 25 51
rect 31 50 35 52
rect 43 51 83 52
rect 31 48 32 50
rect 34 48 35 50
rect 31 47 35 48
rect 21 39 22 41
rect 24 39 25 41
rect 21 37 25 39
rect 28 43 35 47
rect 28 32 32 43
rect 71 38 75 43
rect 71 36 72 38
rect 74 36 75 38
rect 14 31 32 32
rect 14 29 16 31
rect 18 30 32 31
rect 18 29 43 30
rect 14 28 39 29
rect 28 27 39 28
rect 41 27 43 29
rect 28 26 43 27
rect 48 29 52 31
rect 48 27 49 29
rect 51 27 52 29
rect 48 22 52 27
rect 71 34 75 36
rect 79 40 83 51
rect 109 55 113 59
rect 109 51 124 55
rect 79 38 85 40
rect 79 36 82 38
rect 84 36 85 38
rect 79 34 85 36
rect 79 31 83 34
rect 63 27 83 31
rect 63 23 67 27
rect 99 42 105 43
rect 120 38 124 51
rect 127 48 128 59
rect 120 36 121 38
rect 123 36 124 38
rect 120 30 124 36
rect 106 29 124 30
rect 106 27 108 29
rect 110 27 124 29
rect 106 26 124 27
rect 27 21 49 22
rect 18 18 22 20
rect 27 19 29 21
rect 31 20 49 21
rect 51 20 52 22
rect 31 19 52 20
rect 57 22 67 23
rect 57 20 59 22
rect 61 20 67 22
rect 57 19 67 20
rect 27 18 52 19
rect 18 16 19 18
rect 21 16 22 18
rect 96 16 102 17
rect 18 13 22 16
rect 74 15 80 16
rect 74 13 76 15
rect 78 13 80 15
rect 96 14 98 16
rect 100 14 102 16
rect 96 13 102 14
rect 115 16 121 17
rect 115 14 117 16
rect 119 14 121 16
rect 115 13 121 14
rect 26 -5 28 -3
rect 30 -5 32 -3
rect 26 -6 32 -5
rect 84 -6 88 -3
rect 84 -8 85 -6
rect 87 -8 88 -6
rect 54 -9 79 -8
rect 39 -10 49 -9
rect 39 -12 45 -10
rect 47 -12 49 -10
rect 39 -13 49 -12
rect 54 -10 75 -9
rect 54 -12 55 -10
rect 57 -11 75 -10
rect 77 -11 79 -9
rect 84 -10 88 -8
rect 57 -12 79 -11
rect 39 -17 43 -13
rect 23 -21 43 -17
rect 23 -24 27 -21
rect 54 -17 58 -12
rect 54 -19 55 -17
rect 57 -19 58 -17
rect 54 -21 58 -19
rect 63 -17 78 -16
rect 63 -19 65 -17
rect 67 -18 78 -17
rect 67 -19 92 -18
rect 63 -20 88 -19
rect 74 -21 88 -20
rect 90 -21 92 -19
rect 21 -26 27 -24
rect 21 -28 22 -26
rect 24 -28 27 -26
rect 21 -30 27 -28
rect 23 -41 27 -30
rect 31 -26 35 -24
rect 74 -22 92 -21
rect 31 -28 32 -26
rect 34 -28 35 -26
rect 31 -33 35 -28
rect 74 -33 78 -22
rect 71 -37 78 -33
rect 81 -29 85 -27
rect 81 -31 82 -29
rect 84 -31 85 -29
rect 71 -38 75 -37
rect 71 -40 72 -38
rect 74 -40 75 -38
rect 23 -42 63 -41
rect 71 -42 75 -40
rect 81 -41 85 -31
rect 23 -44 37 -42
rect 39 -44 63 -42
rect 23 -45 63 -44
rect 79 -45 85 -41
rect 36 -49 40 -45
rect 59 -49 83 -45
rect 25 -50 31 -49
rect 25 -52 27 -50
rect 29 -52 31 -50
rect 25 -57 31 -52
rect 36 -51 37 -49
rect 39 -51 40 -49
rect 36 -53 40 -51
rect 47 -50 53 -49
rect 47 -52 49 -50
rect 51 -52 53 -50
rect 25 -59 27 -57
rect 29 -59 31 -57
rect 47 -57 53 -52
rect 47 -59 49 -57
rect 51 -59 53 -57
rect 82 -57 88 -56
rect 82 -59 84 -57
rect 86 -59 88 -57
<< via1 >>
rect 8 31 10 33
rect 97 31 99 33
rect 48 -22 50 -20
rect 17 -40 19 -38
<< labels >>
rlabel alu1 53 73 53 73 6 vdd
rlabel alu1 53 9 53 9 1 gnd
rlabel alu1 65 37 65 37 6 a
rlabel alu1 57 45 57 45 1 b
rlabel alu1 97 -27 97 -27 2 so
rlabel alu1 53 -63 53 -63 2 vdd
rlabel alu1 53 1 53 1 5 gnd
rlabel alu1 49 -35 49 -35 1 cin
rlabel alu1 114 73 114 73 4 vdd
rlabel alu1 130 45 130 45 1 co
<< end >>
