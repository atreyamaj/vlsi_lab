magic
tech scmos
timestamp 1553795060
<< ab >>
rect 4 63 181 77
rect 4 59 6 63
rect 8 59 178 63
rect 180 59 181 63
rect 4 5 181 59
rect 183 5 224 77
<< nwell >>
rect -1 37 227 82
<< pwell >>
rect -1 0 227 37
<< poly >>
rect 13 71 15 75
rect 36 68 38 73
rect 43 68 45 73
rect 61 71 63 75
rect 71 71 73 75
rect 81 71 83 75
rect 103 71 105 75
rect 113 71 115 75
rect 123 71 125 75
rect 26 59 28 64
rect 13 33 15 46
rect 26 43 28 46
rect 141 68 143 73
rect 148 68 150 73
rect 171 71 173 75
rect 192 71 194 75
rect 199 71 201 75
rect 158 59 160 64
rect 212 61 214 66
rect 192 47 194 50
rect 158 43 160 46
rect 19 41 28 43
rect 19 39 21 41
rect 23 39 25 41
rect 36 40 38 43
rect 43 40 45 43
rect 61 40 63 43
rect 71 40 73 43
rect 81 40 83 43
rect 103 40 105 43
rect 113 40 115 43
rect 123 40 125 43
rect 141 40 143 43
rect 148 40 150 43
rect 158 41 167 43
rect 19 37 25 39
rect 13 31 19 33
rect 13 29 15 31
rect 17 29 19 31
rect 13 27 19 29
rect 13 24 15 27
rect 23 24 25 37
rect 33 38 39 40
rect 33 36 35 38
rect 37 36 39 38
rect 33 34 39 36
rect 43 38 65 40
rect 43 36 54 38
rect 56 36 61 38
rect 63 36 65 38
rect 43 34 65 36
rect 69 38 75 40
rect 69 36 71 38
rect 73 36 75 38
rect 69 34 75 36
rect 79 38 85 40
rect 79 36 81 38
rect 83 36 85 38
rect 79 34 85 36
rect 101 38 107 40
rect 101 36 103 38
rect 105 36 107 38
rect 101 34 107 36
rect 111 38 117 40
rect 111 36 113 38
rect 115 36 117 38
rect 111 34 117 36
rect 121 38 143 40
rect 121 36 123 38
rect 125 36 130 38
rect 132 36 143 38
rect 121 34 143 36
rect 147 38 153 40
rect 147 36 149 38
rect 151 36 153 38
rect 147 34 153 36
rect 33 31 35 34
rect 43 31 45 34
rect 63 31 65 34
rect 70 31 72 34
rect 13 7 15 11
rect 23 9 25 14
rect 33 12 35 17
rect 43 12 45 17
rect 81 25 83 34
rect 103 25 105 34
rect 114 31 116 34
rect 121 31 123 34
rect 141 31 143 34
rect 151 31 153 34
rect 161 39 163 41
rect 165 39 167 41
rect 161 37 167 39
rect 161 24 163 37
rect 171 33 173 46
rect 188 45 194 47
rect 188 43 190 45
rect 192 43 194 45
rect 188 41 194 43
rect 167 31 173 33
rect 192 31 194 41
rect 199 40 201 50
rect 212 40 214 43
rect 198 38 204 40
rect 198 36 200 38
rect 202 36 204 38
rect 198 34 204 36
rect 208 38 214 40
rect 208 36 210 38
rect 212 36 214 38
rect 208 34 214 36
rect 202 31 204 34
rect 212 31 214 34
rect 167 29 169 31
rect 171 29 173 31
rect 167 27 173 29
rect 171 24 173 27
rect 141 12 143 17
rect 151 12 153 17
rect 63 7 65 11
rect 70 7 72 11
rect 81 7 83 11
rect 103 7 105 11
rect 114 7 116 11
rect 121 7 123 11
rect 161 9 163 14
rect 192 20 194 25
rect 202 20 204 25
rect 212 17 214 22
rect 171 7 173 11
<< ndif >>
rect 28 24 33 31
rect 6 22 13 24
rect 6 20 8 22
rect 10 20 13 22
rect 6 18 13 20
rect 8 11 13 18
rect 15 18 23 24
rect 15 16 18 18
rect 20 16 23 18
rect 15 14 23 16
rect 25 21 33 24
rect 25 19 28 21
rect 30 19 33 21
rect 25 17 33 19
rect 35 29 43 31
rect 35 27 38 29
rect 40 27 43 29
rect 35 17 43 27
rect 45 29 52 31
rect 45 27 48 29
rect 50 27 52 29
rect 45 22 52 27
rect 58 24 63 31
rect 45 20 48 22
rect 50 20 52 22
rect 45 17 52 20
rect 56 22 63 24
rect 56 20 58 22
rect 60 20 63 22
rect 56 18 63 20
rect 25 14 30 17
rect 15 11 20 14
rect 58 11 63 18
rect 65 11 70 31
rect 72 25 79 31
rect 107 25 114 31
rect 72 15 81 25
rect 72 13 75 15
rect 77 13 81 15
rect 72 11 81 13
rect 83 22 90 25
rect 83 20 86 22
rect 88 20 90 22
rect 83 18 90 20
rect 96 22 103 25
rect 96 20 98 22
rect 100 20 103 22
rect 96 18 103 20
rect 83 11 88 18
rect 98 11 103 18
rect 105 15 114 25
rect 105 13 109 15
rect 111 13 114 15
rect 105 11 114 13
rect 116 11 121 31
rect 123 24 128 31
rect 134 29 141 31
rect 134 27 136 29
rect 138 27 141 29
rect 123 22 130 24
rect 123 20 126 22
rect 128 20 130 22
rect 123 18 130 20
rect 134 22 141 27
rect 134 20 136 22
rect 138 20 141 22
rect 123 11 128 18
rect 134 17 141 20
rect 143 29 151 31
rect 143 27 146 29
rect 148 27 151 29
rect 143 17 151 27
rect 153 24 158 31
rect 185 25 192 31
rect 194 29 202 31
rect 194 27 197 29
rect 199 27 202 29
rect 194 25 202 27
rect 204 25 212 31
rect 153 21 161 24
rect 153 19 156 21
rect 158 19 161 21
rect 153 17 161 19
rect 156 14 161 17
rect 163 18 171 24
rect 163 16 166 18
rect 168 16 171 18
rect 163 14 171 16
rect 166 11 171 14
rect 173 22 180 24
rect 173 20 176 22
rect 178 20 180 22
rect 173 18 180 20
rect 185 18 190 25
rect 206 22 212 25
rect 214 29 221 31
rect 214 27 217 29
rect 219 27 221 29
rect 214 25 221 27
rect 214 22 219 25
rect 206 18 210 22
rect 173 11 178 18
rect 185 16 191 18
rect 185 14 187 16
rect 189 14 191 16
rect 185 12 191 14
rect 204 16 210 18
rect 204 14 206 16
rect 208 14 210 16
rect 204 12 210 14
<< pdif >>
rect 8 59 13 71
rect 6 57 13 59
rect 6 55 8 57
rect 10 55 13 57
rect 6 50 13 55
rect 6 48 8 50
rect 10 48 13 50
rect 6 46 13 48
rect 15 69 24 71
rect 15 67 19 69
rect 21 67 24 69
rect 47 69 61 71
rect 47 68 54 69
rect 15 59 24 67
rect 31 59 36 68
rect 15 46 26 59
rect 28 50 36 59
rect 28 48 31 50
rect 33 48 36 50
rect 28 46 36 48
rect 31 43 36 46
rect 38 43 43 68
rect 45 67 54 68
rect 56 67 61 69
rect 45 62 61 67
rect 45 60 54 62
rect 56 60 61 62
rect 45 43 61 60
rect 63 61 71 71
rect 63 59 66 61
rect 68 59 71 61
rect 63 54 71 59
rect 63 52 66 54
rect 68 52 71 54
rect 63 43 71 52
rect 73 69 81 71
rect 73 67 76 69
rect 78 67 81 69
rect 73 62 81 67
rect 73 60 76 62
rect 78 60 81 62
rect 73 43 81 60
rect 83 56 88 71
rect 98 56 103 71
rect 83 54 90 56
rect 83 52 86 54
rect 88 52 90 54
rect 83 47 90 52
rect 83 45 86 47
rect 88 45 90 47
rect 83 43 90 45
rect 96 54 103 56
rect 96 52 98 54
rect 100 52 103 54
rect 96 47 103 52
rect 96 45 98 47
rect 100 45 103 47
rect 96 43 103 45
rect 105 69 113 71
rect 105 67 108 69
rect 110 67 113 69
rect 105 62 113 67
rect 105 60 108 62
rect 110 60 113 62
rect 105 43 113 60
rect 115 61 123 71
rect 115 59 118 61
rect 120 59 123 61
rect 115 54 123 59
rect 115 52 118 54
rect 120 52 123 54
rect 115 43 123 52
rect 125 69 139 71
rect 125 67 130 69
rect 132 68 139 69
rect 162 69 171 71
rect 132 67 141 68
rect 125 62 141 67
rect 125 60 130 62
rect 132 60 141 62
rect 125 43 141 60
rect 143 43 148 68
rect 150 59 155 68
rect 162 67 165 69
rect 167 67 171 69
rect 162 59 171 67
rect 150 50 158 59
rect 150 48 153 50
rect 155 48 158 50
rect 150 46 158 48
rect 160 46 171 59
rect 173 59 178 71
rect 187 64 192 71
rect 185 62 192 64
rect 185 60 187 62
rect 189 60 192 62
rect 173 57 180 59
rect 185 58 192 60
rect 173 55 176 57
rect 178 55 180 57
rect 173 50 180 55
rect 187 50 192 58
rect 194 50 199 71
rect 201 69 210 71
rect 201 67 206 69
rect 208 67 210 69
rect 201 61 210 67
rect 201 50 212 61
rect 173 48 176 50
rect 178 48 180 50
rect 173 46 180 48
rect 150 43 155 46
rect 204 43 212 50
rect 214 59 221 61
rect 214 57 217 59
rect 219 57 221 59
rect 214 52 221 57
rect 214 50 217 52
rect 219 50 221 52
rect 214 48 221 50
rect 214 43 219 48
<< alu1 >>
rect 2 72 224 77
rect 2 70 216 72
rect 218 70 224 72
rect 2 69 224 70
rect 217 63 221 64
rect 208 59 221 63
rect 6 57 11 59
rect 6 55 8 57
rect 10 55 11 57
rect 6 50 11 55
rect 6 48 8 50
rect 10 48 11 50
rect 6 46 11 48
rect 6 30 10 46
rect 37 43 75 47
rect 37 40 42 43
rect 34 38 42 40
rect 34 36 35 38
rect 37 36 42 38
rect 34 34 42 36
rect 52 38 67 39
rect 52 36 54 38
rect 56 36 61 38
rect 63 36 67 38
rect 52 35 67 36
rect 6 28 7 30
rect 9 28 10 30
rect 6 24 10 28
rect 6 22 11 24
rect 54 26 58 35
rect 85 54 91 56
rect 85 52 86 54
rect 88 52 91 54
rect 85 47 91 52
rect 85 45 86 47
rect 88 45 91 47
rect 85 43 91 45
rect 87 38 91 43
rect 87 36 88 38
rect 90 36 91 38
rect 87 23 91 36
rect 6 20 8 22
rect 10 20 11 22
rect 6 18 11 20
rect 85 22 91 23
rect 85 20 86 22
rect 88 20 91 22
rect 85 19 91 20
rect 95 54 101 56
rect 175 57 180 59
rect 175 55 176 57
rect 178 55 180 57
rect 95 52 98 54
rect 100 52 101 54
rect 95 51 101 52
rect 95 49 98 51
rect 100 49 101 51
rect 95 47 101 49
rect 95 45 98 47
rect 100 45 101 47
rect 95 43 101 45
rect 95 23 99 43
rect 111 43 149 47
rect 144 40 149 43
rect 119 38 134 39
rect 119 36 123 38
rect 125 36 130 38
rect 132 36 134 38
rect 119 35 134 36
rect 144 38 152 40
rect 144 36 149 38
rect 151 36 152 38
rect 128 30 132 35
rect 144 34 152 36
rect 175 50 180 55
rect 175 48 176 50
rect 178 48 180 50
rect 175 46 180 48
rect 128 28 129 30
rect 131 28 132 30
rect 128 26 132 28
rect 95 22 101 23
rect 95 20 98 22
rect 100 20 101 22
rect 95 19 101 20
rect 176 24 180 46
rect 185 51 189 56
rect 185 49 186 51
rect 188 49 189 51
rect 185 47 189 49
rect 185 45 206 47
rect 185 43 190 45
rect 192 43 206 45
rect 185 38 206 39
rect 185 36 186 38
rect 188 36 200 38
rect 202 36 206 38
rect 185 35 206 36
rect 219 57 221 59
rect 217 52 221 57
rect 219 50 221 52
rect 185 26 189 35
rect 217 31 221 50
rect 216 29 221 31
rect 216 27 217 29
rect 219 27 221 29
rect 216 25 221 27
rect 175 22 180 24
rect 175 20 176 22
rect 178 20 180 22
rect 175 18 180 20
rect 2 12 224 13
rect 2 10 216 12
rect 218 10 224 12
rect 2 5 224 10
<< alu2 >>
rect 97 51 189 52
rect 97 49 98 51
rect 100 49 186 51
rect 188 49 189 51
rect 97 48 189 49
rect 87 38 190 39
rect 87 36 88 38
rect 90 36 186 38
rect 188 36 190 38
rect 87 35 190 36
rect 6 30 132 31
rect 6 28 7 30
rect 9 28 129 30
rect 131 28 132 30
rect 6 27 132 28
<< ptie >>
rect 214 12 220 14
rect 214 10 216 12
rect 218 10 220 12
rect 214 8 220 10
<< ntie >>
rect 214 72 220 74
rect 214 70 216 72
rect 218 70 220 72
rect 214 68 220 70
<< nmos >>
rect 13 11 15 24
rect 23 14 25 24
rect 33 17 35 31
rect 43 17 45 31
rect 63 11 65 31
rect 70 11 72 31
rect 81 11 83 25
rect 103 11 105 25
rect 114 11 116 31
rect 121 11 123 31
rect 141 17 143 31
rect 151 17 153 31
rect 192 25 194 31
rect 202 25 204 31
rect 161 14 163 24
rect 171 11 173 24
rect 212 22 214 31
<< pmos >>
rect 13 46 15 71
rect 26 46 28 59
rect 36 43 38 68
rect 43 43 45 68
rect 61 43 63 71
rect 71 43 73 71
rect 81 43 83 71
rect 103 43 105 71
rect 113 43 115 71
rect 123 43 125 71
rect 141 43 143 68
rect 148 43 150 68
rect 158 46 160 59
rect 171 46 173 71
rect 192 50 194 71
rect 199 50 201 71
rect 212 43 214 61
<< polyct0 >>
rect 21 39 23 41
rect 15 29 17 31
rect 71 36 73 38
rect 81 36 83 38
rect 103 36 105 38
rect 113 36 115 38
rect 163 39 165 41
rect 210 36 212 38
rect 169 29 171 31
<< polyct1 >>
rect 35 36 37 38
rect 54 36 56 38
rect 61 36 63 38
rect 123 36 125 38
rect 130 36 132 38
rect 149 36 151 38
rect 190 43 192 45
rect 200 36 202 38
<< ndifct0 >>
rect 18 16 20 18
rect 28 19 30 21
rect 38 27 40 29
rect 48 27 50 29
rect 48 20 50 22
rect 58 20 60 22
rect 75 13 77 15
rect 109 13 111 15
rect 136 27 138 29
rect 126 20 128 22
rect 136 20 138 22
rect 146 27 148 29
rect 197 27 199 29
rect 156 19 158 21
rect 166 16 168 18
rect 187 14 189 16
rect 206 14 208 16
<< ndifct1 >>
rect 8 20 10 22
rect 86 20 88 22
rect 98 20 100 22
rect 176 20 178 22
rect 217 27 219 29
<< ntiect1 >>
rect 216 70 218 72
<< ptiect1 >>
rect 216 10 218 12
<< pdifct0 >>
rect 19 67 21 69
rect 31 48 33 50
rect 54 67 56 69
rect 54 60 56 62
rect 66 59 68 61
rect 66 52 68 54
rect 76 67 78 69
rect 76 60 78 62
rect 108 67 110 69
rect 108 60 110 62
rect 118 59 120 61
rect 118 52 120 54
rect 130 67 132 69
rect 130 60 132 62
rect 165 67 167 69
rect 153 48 155 50
rect 187 60 189 62
rect 206 67 208 69
<< pdifct1 >>
rect 8 55 10 57
rect 8 48 10 50
rect 86 52 88 54
rect 86 45 88 47
rect 98 52 100 54
rect 98 45 100 47
rect 176 55 178 57
rect 176 48 178 50
rect 217 57 219 59
rect 217 50 219 52
<< alu0 >>
rect 17 67 19 69
rect 21 67 23 69
rect 17 66 23 67
rect 52 67 54 69
rect 56 67 58 69
rect 52 62 58 67
rect 74 67 76 69
rect 78 67 80 69
rect 52 60 54 62
rect 56 60 58 62
rect 52 59 58 60
rect 65 61 69 63
rect 65 59 66 61
rect 68 59 69 61
rect 74 62 80 67
rect 74 60 76 62
rect 78 60 80 62
rect 74 59 80 60
rect 106 67 108 69
rect 110 67 112 69
rect 106 62 112 67
rect 128 67 130 69
rect 132 67 134 69
rect 106 60 108 62
rect 110 60 112 62
rect 106 59 112 60
rect 117 61 121 63
rect 117 59 118 61
rect 120 59 121 61
rect 128 62 134 67
rect 163 67 165 69
rect 167 67 169 69
rect 163 66 169 67
rect 204 67 206 69
rect 208 67 210 69
rect 204 66 210 67
rect 128 60 130 62
rect 132 60 134 62
rect 128 59 134 60
rect 185 62 202 63
rect 185 60 187 62
rect 189 60 202 62
rect 185 59 202 60
rect 22 55 46 59
rect 65 55 69 59
rect 20 51 26 55
rect 42 54 82 55
rect 42 52 66 54
rect 68 52 82 54
rect 20 41 24 51
rect 30 50 34 52
rect 42 51 82 52
rect 30 48 31 50
rect 33 48 34 50
rect 30 47 34 48
rect 20 39 21 41
rect 23 39 24 41
rect 20 37 24 39
rect 27 43 34 47
rect 27 32 31 43
rect 70 38 74 43
rect 70 36 71 38
rect 73 36 74 38
rect 13 31 31 32
rect 13 29 15 31
rect 17 30 31 31
rect 17 29 42 30
rect 13 28 38 29
rect 27 27 38 28
rect 40 27 42 29
rect 27 26 42 27
rect 47 29 51 31
rect 47 27 48 29
rect 50 27 51 29
rect 47 22 51 27
rect 70 34 74 36
rect 78 40 82 51
rect 78 38 84 40
rect 78 36 81 38
rect 83 36 84 38
rect 78 34 84 36
rect 78 31 82 34
rect 62 27 82 31
rect 62 23 66 27
rect 26 21 48 22
rect 17 18 21 20
rect 26 19 28 21
rect 30 20 48 21
rect 50 20 51 22
rect 30 19 51 20
rect 56 22 66 23
rect 56 20 58 22
rect 60 20 66 22
rect 56 19 66 20
rect 117 55 121 59
rect 140 55 164 59
rect 104 54 144 55
rect 104 52 118 54
rect 120 52 144 54
rect 104 51 144 52
rect 104 40 108 51
rect 152 50 156 52
rect 160 51 166 55
rect 152 48 153 50
rect 155 48 156 50
rect 152 47 156 48
rect 152 43 159 47
rect 102 38 108 40
rect 102 36 103 38
rect 105 36 108 38
rect 102 34 108 36
rect 112 38 116 43
rect 112 36 113 38
rect 115 36 116 38
rect 112 34 116 36
rect 104 31 108 34
rect 104 27 124 31
rect 120 23 124 27
rect 155 32 159 43
rect 162 41 166 51
rect 162 39 163 41
rect 165 39 166 41
rect 162 37 166 39
rect 155 31 173 32
rect 135 29 139 31
rect 155 30 169 31
rect 135 27 136 29
rect 138 27 139 29
rect 120 22 130 23
rect 120 20 126 22
rect 128 20 130 22
rect 120 19 130 20
rect 135 22 139 27
rect 144 29 169 30
rect 171 29 173 31
rect 144 27 146 29
rect 148 28 173 29
rect 148 27 159 28
rect 144 26 159 27
rect 198 55 202 59
rect 198 51 213 55
rect 188 42 194 43
rect 209 38 213 51
rect 216 48 217 59
rect 209 36 210 38
rect 212 36 213 38
rect 209 30 213 36
rect 195 29 213 30
rect 195 27 197 29
rect 199 27 213 29
rect 195 26 213 27
rect 135 20 136 22
rect 138 21 160 22
rect 138 20 156 21
rect 135 19 156 20
rect 158 19 160 21
rect 26 18 51 19
rect 135 18 160 19
rect 165 18 169 20
rect 17 16 18 18
rect 20 16 21 18
rect 165 16 166 18
rect 168 16 169 18
rect 17 13 21 16
rect 73 15 79 16
rect 73 13 75 15
rect 77 13 79 15
rect 107 15 113 16
rect 107 13 109 15
rect 111 13 113 15
rect 165 13 169 16
rect 185 16 191 17
rect 185 14 187 16
rect 189 14 191 16
rect 185 13 191 14
rect 204 16 210 17
rect 204 14 206 16
rect 208 14 210 16
rect 204 13 210 14
<< via1 >>
rect 7 28 9 30
rect 88 36 90 38
rect 98 49 100 51
rect 129 28 131 30
rect 186 49 188 51
rect 186 36 188 38
<< labels >>
rlabel alu1 52 73 52 73 6 vdd
rlabel alu1 52 9 52 9 1 gnd
rlabel alu1 64 37 64 37 6 a
rlabel alu1 56 45 56 45 1 b
rlabel alu1 134 9 134 9 1 gnd
rlabel alu1 134 73 134 73 4 vdd
rlabel alu1 178 37 178 37 4 so
rlabel alu1 131 45 131 45 1 cin
rlabel alu1 203 73 203 73 4 vdd
rlabel alu1 219 43 219 43 1 cout
<< end >>
