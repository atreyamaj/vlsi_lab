* Inverter using a NMOS Transistor

.include ./t14y_tsmc_025_level3.txt

* NET List
* m0 drain gate source bulk
m0 out in 0 0 cmosn l=2.5u w=10u
rl supply out 7k
cl out 0 5n

* source
vdd supply 0 dc 3.3
vin in 0 dc 3.3 pulse(0 3.3 0 0.1n 0.1n 0.5m 1m)

.control

dc vin 0 3.3 0.01
plot out

plot deriv(out)
meas dc vol find out when in=3.29
let slope=deriv(out)
let voh=3.3
meas dc vih find in when slope=-1 cross=2
meas dc vil find in when slope=-1 cross=1

let v90 = voh-0.1*(voh-vol)
let v10 = vol+0.1*(voh-vol)
let vhalf = voh-0.5*(voh-vol)

tran 0.1m 4m
plot in out
plot -vdd#branch
meas tran trise trig out val=dc1.v10 rise=1 targ out val=dc1.v90 rise=1
meas tran tfall trig out val=dc1.v90 fall=1 targ out val=dc1.v10 fall=1

meas tran thl trig out val=dc1.vhalf rise=1 targ out val=dc1.vhalf fall=2
meas tran tlh trig out val=dc1.vhalf fall=1 targ out val=dc1.vhalf rise=1
let td = 0.5*(thl+tlh)

let power = -3.3*vdd#branch
meas tran pavg AVG power from=0m to=2m 

.endc
.end
